magic
tech sky130A
magscale 1 2
timestamp 1654931914
<< metal1 >>
rect 3878 700748 3884 700800
rect 3936 700788 3942 700800
rect 8110 700788 8116 700800
rect 3936 700760 8116 700788
rect 3936 700748 3942 700760
rect 8110 700748 8116 700760
rect 8168 700748 8174 700800
rect 102042 700748 102048 700800
rect 102100 700788 102106 700800
rect 105446 700788 105452 700800
rect 102100 700760 105452 700788
rect 102100 700748 102106 700760
rect 105446 700748 105452 700760
rect 105504 700748 105510 700800
rect 200022 700748 200028 700800
rect 200080 700788 200086 700800
rect 202782 700788 202788 700800
rect 200080 700760 202788 700788
rect 200080 700748 200086 700760
rect 202782 700748 202788 700760
rect 202840 700748 202846 700800
rect 314470 700748 314476 700800
rect 314528 700788 314534 700800
rect 316310 700788 316316 700800
rect 314528 700760 316316 700788
rect 314528 700748 314534 700760
rect 316310 700748 316316 700760
rect 316368 700748 316374 700800
rect 363506 700408 363512 700460
rect 363564 700448 363570 700460
rect 364978 700448 364984 700460
rect 363564 700420 364984 700448
rect 363564 700408 363570 700420
rect 364978 700408 364984 700420
rect 365036 700408 365042 700460
rect 412450 700408 412456 700460
rect 412508 700448 412514 700460
rect 413646 700448 413652 700460
rect 412508 700420 413652 700448
rect 412508 700408 412514 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 20346 700204 20352 700256
rect 20404 700244 20410 700256
rect 24302 700244 24308 700256
rect 20404 700216 24308 700244
rect 20404 700204 20410 700216
rect 24302 700204 24308 700216
rect 24360 700204 24366 700256
rect 36722 700204 36728 700256
rect 36780 700244 36786 700256
rect 40494 700244 40500 700256
rect 36780 700216 40500 700244
rect 36780 700204 36786 700216
rect 40494 700204 40500 700216
rect 40552 700204 40558 700256
rect 69382 700204 69388 700256
rect 69440 700244 69446 700256
rect 72970 700244 72976 700256
rect 69440 700216 72976 700244
rect 69440 700204 69446 700216
rect 72970 700204 72976 700216
rect 73028 700204 73034 700256
rect 85758 700204 85764 700256
rect 85816 700244 85822 700256
rect 89162 700244 89168 700256
rect 85816 700216 89168 700244
rect 85816 700204 85822 700216
rect 89162 700204 89168 700216
rect 89220 700204 89226 700256
rect 134702 700204 134708 700256
rect 134760 700244 134766 700256
rect 137830 700244 137836 700256
rect 134760 700216 137836 700244
rect 134760 700204 134766 700216
rect 137830 700204 137836 700216
rect 137888 700204 137894 700256
rect 167362 700204 167368 700256
rect 167420 700244 167426 700256
rect 170306 700244 170312 700256
rect 167420 700216 170312 700244
rect 167420 700204 167426 700216
rect 170306 700204 170312 700216
rect 170364 700204 170370 700256
rect 183738 700204 183744 700256
rect 183796 700244 183802 700256
rect 186498 700244 186504 700256
rect 183796 700216 186504 700244
rect 183796 700204 183802 700216
rect 186498 700204 186504 700216
rect 186556 700204 186562 700256
rect 232774 700204 232780 700256
rect 232832 700244 232838 700256
rect 235166 700244 235172 700256
rect 232832 700216 235172 700244
rect 232832 700204 232838 700216
rect 235166 700204 235172 700216
rect 235224 700204 235230 700256
rect 249058 700204 249064 700256
rect 249116 700244 249122 700256
rect 251450 700244 251456 700256
rect 249116 700216 251456 700244
rect 249116 700204 249122 700216
rect 251450 700204 251456 700216
rect 251508 700204 251514 700256
rect 265434 700204 265440 700256
rect 265492 700244 265498 700256
rect 267642 700244 267648 700256
rect 265492 700216 267648 700244
rect 265492 700204 265498 700216
rect 267642 700204 267648 700216
rect 267700 700204 267706 700256
rect 281810 700204 281816 700256
rect 281868 700244 281874 700256
rect 283834 700244 283840 700256
rect 281868 700216 283840 700244
rect 281868 700204 281874 700216
rect 283834 700204 283840 700216
rect 283892 700204 283898 700256
rect 330754 700204 330760 700256
rect 330812 700244 330818 700256
rect 332502 700244 332508 700256
rect 330812 700216 332508 700244
rect 330812 700204 330818 700216
rect 332502 700204 332508 700216
rect 332560 700204 332566 700256
rect 347130 700204 347136 700256
rect 347188 700244 347194 700256
rect 348786 700244 348792 700256
rect 347188 700216 348792 700244
rect 347188 700204 347194 700216
rect 348786 700204 348792 700216
rect 348844 700204 348850 700256
rect 396166 700204 396172 700256
rect 396224 700244 396230 700256
rect 397454 700244 397460 700256
rect 396224 700216 397460 700244
rect 396224 700204 396230 700216
rect 397454 700204 397460 700216
rect 397512 700204 397518 700256
rect 428826 700204 428832 700256
rect 428884 700244 428890 700256
rect 429838 700244 429844 700256
rect 428884 700216 429844 700244
rect 428884 700204 428890 700216
rect 429838 700204 429844 700216
rect 429896 700204 429902 700256
rect 445202 700204 445208 700256
rect 445260 700244 445266 700256
rect 446122 700244 446128 700256
rect 445260 700216 446128 700244
rect 445260 700204 445266 700216
rect 446122 700204 446128 700216
rect 446180 700204 446186 700256
rect 461486 700204 461492 700256
rect 461544 700244 461550 700256
rect 462314 700244 462320 700256
rect 461544 700216 462320 700244
rect 461544 700204 461550 700216
rect 462314 700204 462320 700216
rect 462372 700204 462378 700256
rect 118418 700136 118424 700188
rect 118476 700176 118482 700188
rect 121638 700176 121644 700188
rect 118476 700148 121644 700176
rect 118476 700136 118482 700148
rect 121638 700136 121644 700148
rect 121696 700136 121702 700188
rect 151078 700136 151084 700188
rect 151136 700176 151142 700188
rect 154114 700176 154120 700188
rect 151136 700148 154120 700176
rect 151136 700136 151142 700148
rect 154114 700136 154120 700148
rect 154172 700136 154178 700188
rect 216398 700136 216404 700188
rect 216456 700176 216462 700188
rect 218974 700176 218980 700188
rect 216456 700148 218980 700176
rect 216456 700136 216462 700148
rect 218974 700136 218980 700148
rect 219032 700136 219038 700188
rect 298002 700136 298008 700188
rect 298060 700176 298066 700188
rect 300118 700176 300124 700188
rect 298060 700148 300124 700176
rect 298060 700136 298066 700148
rect 300118 700136 300124 700148
rect 300176 700136 300182 700188
rect 477862 700136 477868 700188
rect 477920 700176 477926 700188
rect 478506 700176 478512 700188
rect 477920 700148 478512 700176
rect 477920 700136 477926 700148
rect 478506 700136 478512 700148
rect 478564 700136 478570 700188
rect 494238 700136 494244 700188
rect 494296 700176 494302 700188
rect 494790 700176 494796 700188
rect 494296 700148 494796 700176
rect 494296 700136 494302 700148
rect 494790 700136 494796 700148
rect 494848 700136 494854 700188
rect 53006 700000 53012 700052
rect 53064 700040 53070 700052
rect 56778 700040 56784 700052
rect 53064 700012 56784 700040
rect 53064 700000 53070 700012
rect 56778 700000 56784 700012
rect 56836 700000 56842 700052
rect 379790 699864 379796 699916
rect 379848 699904 379854 699916
rect 381170 699904 381176 699916
rect 379848 699876 381176 699904
rect 379848 699864 379854 699876
rect 381170 699864 381176 699876
rect 381228 699864 381234 699916
rect 578326 644512 578332 644564
rect 578384 644552 578390 644564
rect 580902 644552 580908 644564
rect 578384 644524 580908 644552
rect 578384 644512 578390 644524
rect 580902 644512 580908 644524
rect 580960 644512 580966 644564
rect 578878 257796 578884 257848
rect 578936 257836 578942 257848
rect 580902 257836 580908 257848
rect 578936 257808 580908 257836
rect 578936 257796 578942 257808
rect 580902 257796 580908 257808
rect 580960 257796 580966 257848
rect 578510 151444 578516 151496
rect 578568 151484 578574 151496
rect 580902 151484 580908 151496
rect 578568 151456 580908 151484
rect 578568 151444 578574 151456
rect 580902 151444 580908 151456
rect 580960 151444 580966 151496
rect 578326 44956 578332 45008
rect 578384 44996 578390 45008
rect 579982 44996 579988 45008
rect 578384 44968 579988 44996
rect 578384 44956 578390 44968
rect 579982 44956 579988 44968
rect 580040 44956 580046 45008
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 14502 3924 14508 3936
rect 11204 3896 14508 3924
rect 11204 3884 11210 3896
rect 14502 3884 14508 3896
rect 14560 3884 14566 3936
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 17998 3924 18004 3936
rect 14792 3896 18004 3924
rect 14792 3884 14798 3896
rect 17998 3884 18004 3896
rect 18056 3884 18062 3936
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 23794 3924 23800 3936
rect 20680 3896 23800 3924
rect 20680 3884 20686 3896
rect 23794 3884 23800 3896
rect 23852 3884 23858 3936
rect 24210 3884 24216 3936
rect 24268 3924 24274 3936
rect 27290 3924 27296 3936
rect 24268 3896 27296 3924
rect 24268 3884 24274 3896
rect 27290 3884 27296 3896
rect 27348 3884 27354 3936
rect 27706 3884 27712 3936
rect 27764 3924 27770 3936
rect 30694 3924 30700 3936
rect 27764 3896 30700 3924
rect 27764 3884 27770 3896
rect 30694 3884 30700 3896
rect 30752 3884 30758 3936
rect 32398 3884 32404 3936
rect 32456 3924 32462 3936
rect 35386 3924 35392 3936
rect 32456 3896 35392 3924
rect 32456 3884 32462 3896
rect 35386 3884 35392 3896
rect 35444 3884 35450 3936
rect 38378 3884 38384 3936
rect 38436 3924 38442 3936
rect 41182 3924 41188 3936
rect 38436 3896 41188 3924
rect 38436 3884 38442 3896
rect 41182 3884 41188 3896
rect 41240 3884 41246 3936
rect 43070 3884 43076 3936
rect 43128 3924 43134 3936
rect 45782 3924 45788 3936
rect 43128 3896 45788 3924
rect 43128 3884 43134 3896
rect 45782 3884 45788 3896
rect 45840 3884 45846 3936
rect 46658 3884 46664 3936
rect 46716 3924 46722 3936
rect 49278 3924 49284 3936
rect 46716 3896 49284 3924
rect 46716 3884 46722 3896
rect 49278 3884 49284 3896
rect 49336 3884 49342 3936
rect 50154 3884 50160 3936
rect 50212 3924 50218 3936
rect 52774 3924 52780 3936
rect 50212 3896 52780 3924
rect 50212 3884 50218 3896
rect 52774 3884 52780 3896
rect 52832 3884 52838 3936
rect 56042 3884 56048 3936
rect 56100 3924 56106 3936
rect 58570 3924 58576 3936
rect 56100 3896 58576 3924
rect 56100 3884 56106 3896
rect 58570 3884 58576 3896
rect 58628 3884 58634 3936
rect 72602 3884 72608 3936
rect 72660 3924 72666 3936
rect 74854 3924 74860 3936
rect 72660 3896 74860 3924
rect 72660 3884 72666 3896
rect 74854 3884 74860 3896
rect 74912 3884 74918 3936
rect 247630 3884 247636 3936
rect 247688 3924 247694 3936
rect 248598 3924 248604 3936
rect 247688 3896 248604 3924
rect 247688 3884 247694 3896
rect 248598 3884 248604 3896
rect 248656 3884 248662 3936
rect 285902 3884 285908 3936
rect 285960 3924 285966 3936
rect 287790 3924 287796 3936
rect 285960 3896 287796 3924
rect 285960 3884 285966 3896
rect 287790 3884 287796 3896
rect 287848 3884 287854 3936
rect 1670 3816 1676 3868
rect 1728 3856 1734 3868
rect 5210 3856 5216 3868
rect 1728 3828 5216 3856
rect 1728 3816 1734 3828
rect 5210 3816 5216 3828
rect 5268 3816 5274 3868
rect 13538 3816 13544 3868
rect 13596 3856 13602 3868
rect 16802 3856 16808 3868
rect 13596 3828 16808 3856
rect 13596 3816 13602 3828
rect 16802 3816 16808 3828
rect 16860 3816 16866 3868
rect 19426 3816 19432 3868
rect 19484 3856 19490 3868
rect 22598 3856 22604 3868
rect 19484 3828 22604 3856
rect 19484 3816 19490 3828
rect 22598 3816 22604 3828
rect 22656 3816 22662 3868
rect 23014 3816 23020 3868
rect 23072 3856 23078 3868
rect 26094 3856 26100 3868
rect 23072 3828 26100 3856
rect 23072 3816 23078 3828
rect 26094 3816 26100 3828
rect 26152 3816 26158 3868
rect 26510 3816 26516 3868
rect 26568 3856 26574 3868
rect 29590 3856 29596 3868
rect 26568 3828 29596 3856
rect 26568 3816 26574 3828
rect 29590 3816 29596 3828
rect 29648 3816 29654 3868
rect 30098 3816 30104 3868
rect 30156 3856 30162 3868
rect 33086 3856 33092 3868
rect 30156 3828 33092 3856
rect 30156 3816 30162 3828
rect 33086 3816 33092 3828
rect 33144 3816 33150 3868
rect 33594 3816 33600 3868
rect 33652 3856 33658 3868
rect 36582 3856 36588 3868
rect 33652 3828 36588 3856
rect 33652 3816 33658 3828
rect 36582 3816 36588 3828
rect 36640 3816 36646 3868
rect 37182 3816 37188 3868
rect 37240 3856 37246 3868
rect 39986 3856 39992 3868
rect 37240 3828 39992 3856
rect 37240 3816 37246 3828
rect 39986 3816 39992 3828
rect 40044 3816 40050 3868
rect 41874 3816 41880 3868
rect 41932 3856 41938 3868
rect 44678 3856 44684 3868
rect 41932 3828 44684 3856
rect 41932 3816 41938 3828
rect 44678 3816 44684 3828
rect 44736 3816 44742 3868
rect 45462 3816 45468 3868
rect 45520 3856 45526 3868
rect 48174 3856 48180 3868
rect 45520 3828 48180 3856
rect 45520 3816 45526 3828
rect 48174 3816 48180 3828
rect 48232 3816 48238 3868
rect 48958 3816 48964 3868
rect 49016 3856 49022 3868
rect 51578 3856 51584 3868
rect 49016 3828 51584 3856
rect 49016 3816 49022 3828
rect 51578 3816 51584 3828
rect 51636 3816 51642 3868
rect 53742 3816 53748 3868
rect 53800 3856 53806 3868
rect 56270 3856 56276 3868
rect 53800 3828 56276 3856
rect 53800 3816 53806 3828
rect 56270 3816 56276 3828
rect 56328 3816 56334 3868
rect 57238 3816 57244 3868
rect 57296 3856 57302 3868
rect 59766 3856 59772 3868
rect 57296 3828 59772 3856
rect 57296 3816 57302 3828
rect 59766 3816 59772 3828
rect 59824 3816 59830 3868
rect 71498 3816 71504 3868
rect 71556 3856 71562 3868
rect 73658 3856 73664 3868
rect 71556 3828 73664 3856
rect 71556 3816 71562 3828
rect 73658 3816 73664 3828
rect 73716 3816 73722 3868
rect 78582 3816 78588 3868
rect 78640 3856 78646 3868
rect 80650 3856 80656 3868
rect 78640 3828 80656 3856
rect 78640 3816 78646 3828
rect 80650 3816 80656 3828
rect 80708 3816 80714 3868
rect 80882 3816 80888 3868
rect 80940 3856 80946 3868
rect 82950 3856 82956 3868
rect 80940 3828 82956 3856
rect 80940 3816 80946 3828
rect 82950 3816 82956 3828
rect 83008 3816 83014 3868
rect 87966 3816 87972 3868
rect 88024 3856 88030 3868
rect 89942 3856 89948 3868
rect 88024 3828 89948 3856
rect 88024 3816 88030 3828
rect 89942 3816 89948 3828
rect 90000 3816 90006 3868
rect 96246 3816 96252 3868
rect 96304 3856 96310 3868
rect 98038 3856 98044 3868
rect 96304 3828 98044 3856
rect 96304 3816 96310 3828
rect 98038 3816 98044 3828
rect 98096 3816 98102 3868
rect 244134 3816 244140 3868
rect 244192 3856 244198 3868
rect 245194 3856 245200 3868
rect 244192 3828 245200 3856
rect 244192 3816 244198 3828
rect 245194 3816 245200 3828
rect 245252 3816 245258 3868
rect 256922 3816 256928 3868
rect 256980 3856 256986 3868
rect 258258 3856 258264 3868
rect 256980 3828 258264 3856
rect 256980 3816 256986 3828
rect 258258 3816 258264 3828
rect 258316 3816 258322 3868
rect 259222 3816 259228 3868
rect 259280 3856 259286 3868
rect 260650 3856 260656 3868
rect 259280 3828 260656 3856
rect 259280 3816 259286 3828
rect 260650 3816 260656 3828
rect 260708 3816 260714 3868
rect 261614 3816 261620 3868
rect 261672 3856 261678 3868
rect 262950 3856 262956 3868
rect 261672 3828 262956 3856
rect 261672 3816 261678 3828
rect 262950 3816 262956 3828
rect 263008 3816 263014 3868
rect 263914 3816 263920 3868
rect 263972 3856 263978 3868
rect 265342 3856 265348 3868
rect 263972 3828 265348 3856
rect 263972 3816 263978 3828
rect 265342 3816 265348 3828
rect 265400 3816 265406 3868
rect 268514 3816 268520 3868
rect 268572 3856 268578 3868
rect 270034 3856 270040 3868
rect 268572 3828 270040 3856
rect 268572 3816 268578 3828
rect 270034 3816 270040 3828
rect 270092 3816 270098 3868
rect 270814 3816 270820 3868
rect 270872 3856 270878 3868
rect 272426 3856 272432 3868
rect 270872 3828 272432 3856
rect 270872 3816 270878 3828
rect 272426 3816 272432 3828
rect 272484 3816 272490 3868
rect 275506 3816 275512 3868
rect 275564 3856 275570 3868
rect 277118 3856 277124 3868
rect 275564 3828 277124 3856
rect 275564 3816 275570 3828
rect 277118 3816 277124 3828
rect 277176 3816 277182 3868
rect 277806 3816 277812 3868
rect 277864 3856 277870 3868
rect 279510 3856 279516 3868
rect 277864 3828 279516 3856
rect 277864 3816 277870 3828
rect 279510 3816 279516 3828
rect 279568 3816 279574 3868
rect 284798 3816 284804 3868
rect 284856 3856 284862 3868
rect 286594 3856 286600 3868
rect 284856 3828 286600 3856
rect 284856 3816 284862 3828
rect 286594 3816 286600 3828
rect 286652 3816 286658 3868
rect 292894 3816 292900 3868
rect 292952 3856 292958 3868
rect 294874 3856 294880 3868
rect 292952 3828 294880 3856
rect 292952 3816 292958 3828
rect 294874 3816 294880 3828
rect 294932 3816 294938 3868
rect 299886 3816 299892 3868
rect 299944 3856 299950 3868
rect 301958 3856 301964 3868
rect 299944 3828 301964 3856
rect 299944 3816 299950 3828
rect 301958 3816 301964 3828
rect 302016 3816 302022 3868
rect 306786 3816 306792 3868
rect 306844 3856 306850 3868
rect 309042 3856 309048 3868
rect 306844 3828 309048 3856
rect 306844 3816 306850 3828
rect 309042 3816 309048 3828
rect 309100 3816 309106 3868
rect 566 3748 572 3800
rect 624 3788 630 3800
rect 4106 3788 4112 3800
rect 624 3760 4112 3788
rect 624 3748 630 3760
rect 4106 3748 4112 3760
rect 4164 3748 4170 3800
rect 7650 3748 7656 3800
rect 7708 3788 7714 3800
rect 11006 3788 11012 3800
rect 7708 3760 11012 3788
rect 7708 3748 7714 3760
rect 11006 3748 11012 3760
rect 11064 3748 11070 3800
rect 12342 3748 12348 3800
rect 12400 3788 12406 3800
rect 15698 3788 15704 3800
rect 12400 3760 15704 3788
rect 12400 3748 12406 3760
rect 15698 3748 15704 3760
rect 15756 3748 15762 3800
rect 15930 3748 15936 3800
rect 15988 3788 15994 3800
rect 19102 3788 19108 3800
rect 15988 3760 19108 3788
rect 15988 3748 15994 3760
rect 19102 3748 19108 3760
rect 19160 3748 19166 3800
rect 21818 3748 21824 3800
rect 21876 3788 21882 3800
rect 24898 3788 24904 3800
rect 21876 3760 24904 3788
rect 21876 3748 21882 3760
rect 24898 3748 24904 3760
rect 24956 3748 24962 3800
rect 25314 3748 25320 3800
rect 25372 3788 25378 3800
rect 28394 3788 28400 3800
rect 25372 3760 28400 3788
rect 25372 3748 25378 3760
rect 28394 3748 28400 3760
rect 28452 3748 28458 3800
rect 31294 3748 31300 3800
rect 31352 3788 31358 3800
rect 34190 3788 34196 3800
rect 31352 3760 34196 3788
rect 31352 3748 31358 3760
rect 34190 3748 34196 3760
rect 34248 3748 34254 3800
rect 34790 3748 34796 3800
rect 34848 3788 34854 3800
rect 37686 3788 37692 3800
rect 34848 3760 37692 3788
rect 34848 3748 34854 3760
rect 37686 3748 37692 3760
rect 37744 3748 37750 3800
rect 40678 3748 40684 3800
rect 40736 3788 40742 3800
rect 43482 3788 43488 3800
rect 40736 3760 43488 3788
rect 40736 3748 40742 3760
rect 43482 3748 43488 3760
rect 43540 3748 43546 3800
rect 44266 3748 44272 3800
rect 44324 3788 44330 3800
rect 46978 3788 46984 3800
rect 44324 3760 46984 3788
rect 44324 3748 44330 3760
rect 46978 3748 46984 3760
rect 47036 3748 47042 3800
rect 47854 3748 47860 3800
rect 47912 3788 47918 3800
rect 50474 3788 50480 3800
rect 47912 3760 50480 3788
rect 47912 3748 47918 3760
rect 50474 3748 50480 3760
rect 50532 3748 50538 3800
rect 51350 3748 51356 3800
rect 51408 3788 51414 3800
rect 53970 3788 53976 3800
rect 51408 3760 53976 3788
rect 51408 3748 51414 3760
rect 53970 3748 53976 3760
rect 54028 3748 54034 3800
rect 54938 3748 54944 3800
rect 54996 3788 55002 3800
rect 57374 3788 57380 3800
rect 54996 3760 57380 3788
rect 54996 3748 55002 3760
rect 57374 3748 57380 3760
rect 57432 3748 57438 3800
rect 58434 3748 58440 3800
rect 58492 3788 58498 3800
rect 60870 3788 60876 3800
rect 58492 3760 60876 3788
rect 58492 3748 58498 3760
rect 60870 3748 60876 3760
rect 60928 3748 60934 3800
rect 64322 3748 64328 3800
rect 64380 3788 64386 3800
rect 66666 3788 66672 3800
rect 64380 3760 66672 3788
rect 64380 3748 64386 3760
rect 66666 3748 66672 3760
rect 66724 3748 66730 3800
rect 67082 3748 67088 3800
rect 67140 3788 67146 3800
rect 69058 3788 69064 3800
rect 67140 3760 69064 3788
rect 67140 3748 67146 3760
rect 69058 3748 69064 3760
rect 69116 3748 69122 3800
rect 70302 3748 70308 3800
rect 70360 3788 70366 3800
rect 72462 3788 72468 3800
rect 70360 3760 72468 3788
rect 70360 3748 70366 3760
rect 72462 3748 72468 3760
rect 72520 3748 72526 3800
rect 73798 3748 73804 3800
rect 73856 3788 73862 3800
rect 75958 3788 75964 3800
rect 73856 3760 75964 3788
rect 73856 3748 73862 3760
rect 75958 3748 75964 3760
rect 76016 3748 76022 3800
rect 79686 3748 79692 3800
rect 79744 3788 79750 3800
rect 81754 3788 81760 3800
rect 79744 3760 81760 3788
rect 79744 3748 79750 3760
rect 81754 3748 81760 3760
rect 81812 3748 81818 3800
rect 86862 3748 86868 3800
rect 86920 3788 86926 3800
rect 88746 3788 88752 3800
rect 86920 3760 88752 3788
rect 86920 3748 86926 3760
rect 88746 3748 88752 3760
rect 88804 3748 88810 3800
rect 95142 3748 95148 3800
rect 95200 3788 95206 3800
rect 96842 3788 96848 3800
rect 95200 3760 96848 3788
rect 95200 3748 95206 3760
rect 96842 3748 96848 3760
rect 96900 3748 96906 3800
rect 103330 3748 103336 3800
rect 103388 3788 103394 3800
rect 104938 3788 104944 3800
rect 103388 3760 104944 3788
rect 103388 3748 103394 3760
rect 104938 3748 104944 3760
rect 104996 3748 105002 3800
rect 216350 3748 216356 3800
rect 216408 3788 216414 3800
rect 216858 3788 216864 3800
rect 216408 3760 216864 3788
rect 216408 3748 216414 3760
rect 216858 3748 216864 3760
rect 216916 3748 216922 3800
rect 222146 3748 222152 3800
rect 222204 3788 222210 3800
rect 222746 3788 222752 3800
rect 222204 3760 222752 3788
rect 222204 3748 222210 3760
rect 222746 3748 222752 3760
rect 222804 3748 222810 3800
rect 224446 3748 224452 3800
rect 224504 3788 224510 3800
rect 225138 3788 225144 3800
rect 224504 3760 225144 3788
rect 224504 3748 224510 3760
rect 225138 3748 225144 3760
rect 225196 3748 225202 3800
rect 230242 3748 230248 3800
rect 230300 3788 230306 3800
rect 231026 3788 231032 3800
rect 230300 3760 231032 3788
rect 230300 3748 230306 3760
rect 231026 3748 231032 3760
rect 231084 3748 231090 3800
rect 231438 3748 231444 3800
rect 231496 3788 231502 3800
rect 232222 3788 232228 3800
rect 231496 3760 232228 3788
rect 231496 3748 231502 3760
rect 232222 3748 232228 3760
rect 232280 3748 232286 3800
rect 232542 3748 232548 3800
rect 232600 3788 232606 3800
rect 233418 3788 233424 3800
rect 232600 3760 233424 3788
rect 232600 3748 232606 3760
rect 233418 3748 233424 3760
rect 233476 3748 233482 3800
rect 233738 3748 233744 3800
rect 233796 3788 233802 3800
rect 234614 3788 234620 3800
rect 233796 3760 234620 3788
rect 233796 3748 233802 3760
rect 234614 3748 234620 3760
rect 234672 3748 234678 3800
rect 237234 3748 237240 3800
rect 237292 3788 237298 3800
rect 238110 3788 238116 3800
rect 237292 3760 238116 3788
rect 237292 3748 237298 3760
rect 238110 3748 238116 3760
rect 238168 3748 238174 3800
rect 238338 3748 238344 3800
rect 238396 3788 238402 3800
rect 239306 3788 239312 3800
rect 238396 3760 239312 3788
rect 238396 3748 238402 3760
rect 239306 3748 239312 3760
rect 239364 3748 239370 3800
rect 239534 3748 239540 3800
rect 239592 3788 239598 3800
rect 240502 3788 240508 3800
rect 239592 3760 240508 3788
rect 239592 3748 239598 3760
rect 240502 3748 240508 3760
rect 240560 3748 240566 3800
rect 240730 3748 240736 3800
rect 240788 3788 240794 3800
rect 241698 3788 241704 3800
rect 240788 3760 241704 3788
rect 240788 3748 240794 3760
rect 241698 3748 241704 3760
rect 241756 3748 241762 3800
rect 241834 3748 241840 3800
rect 241892 3788 241898 3800
rect 242894 3788 242900 3800
rect 241892 3760 242900 3788
rect 241892 3748 241898 3760
rect 242894 3748 242900 3760
rect 242952 3748 242958 3800
rect 245330 3748 245336 3800
rect 245388 3788 245394 3800
rect 246390 3788 246396 3800
rect 245388 3760 246396 3788
rect 245388 3748 245394 3760
rect 246390 3748 246396 3760
rect 246448 3748 246454 3800
rect 246526 3748 246532 3800
rect 246584 3788 246590 3800
rect 247586 3788 247592 3800
rect 246584 3760 247592 3788
rect 246584 3748 246590 3760
rect 247586 3748 247592 3760
rect 247644 3748 247650 3800
rect 250022 3748 250028 3800
rect 250080 3788 250086 3800
rect 251174 3788 251180 3800
rect 250080 3760 251180 3788
rect 250080 3748 250086 3760
rect 251174 3748 251180 3760
rect 251232 3748 251238 3800
rect 252322 3748 252328 3800
rect 252380 3788 252386 3800
rect 253474 3788 253480 3800
rect 252380 3760 253480 3788
rect 252380 3748 252386 3760
rect 253474 3748 253480 3760
rect 253532 3748 253538 3800
rect 255818 3748 255824 3800
rect 255876 3788 255882 3800
rect 257062 3788 257068 3800
rect 255876 3760 257068 3788
rect 255876 3748 255882 3760
rect 257062 3748 257068 3760
rect 257120 3748 257126 3800
rect 258118 3748 258124 3800
rect 258176 3788 258182 3800
rect 259454 3788 259460 3800
rect 258176 3760 259460 3788
rect 258176 3748 258182 3760
rect 259454 3748 259460 3760
rect 259512 3748 259518 3800
rect 260418 3748 260424 3800
rect 260476 3788 260482 3800
rect 261754 3788 261760 3800
rect 260476 3760 261760 3788
rect 260476 3748 260482 3760
rect 261754 3748 261760 3760
rect 261812 3748 261818 3800
rect 262718 3748 262724 3800
rect 262776 3788 262782 3800
rect 264146 3788 264152 3800
rect 262776 3760 264152 3788
rect 262776 3748 262782 3760
rect 264146 3748 264152 3760
rect 264204 3748 264210 3800
rect 265018 3748 265024 3800
rect 265076 3788 265082 3800
rect 266538 3788 266544 3800
rect 265076 3760 266544 3788
rect 265076 3748 265082 3760
rect 266538 3748 266544 3760
rect 266596 3748 266602 3800
rect 267410 3748 267416 3800
rect 267468 3788 267474 3800
rect 268838 3788 268844 3800
rect 267468 3760 268844 3788
rect 267468 3748 267474 3760
rect 268838 3748 268844 3760
rect 268896 3748 268902 3800
rect 269710 3748 269716 3800
rect 269768 3788 269774 3800
rect 271230 3788 271236 3800
rect 269768 3760 271236 3788
rect 269768 3748 269774 3760
rect 271230 3748 271236 3760
rect 271288 3748 271294 3800
rect 272010 3748 272016 3800
rect 272068 3788 272074 3800
rect 273622 3788 273628 3800
rect 272068 3760 273628 3788
rect 272068 3748 272074 3760
rect 273622 3748 273628 3760
rect 273680 3748 273686 3800
rect 276702 3748 276708 3800
rect 276760 3788 276766 3800
rect 278314 3788 278320 3800
rect 276760 3760 278320 3788
rect 276760 3748 276766 3760
rect 278314 3748 278320 3760
rect 278372 3748 278378 3800
rect 279002 3748 279008 3800
rect 279060 3788 279066 3800
rect 280706 3788 280712 3800
rect 279060 3760 280712 3788
rect 279060 3748 279066 3760
rect 280706 3748 280712 3760
rect 280764 3748 280770 3800
rect 283602 3748 283608 3800
rect 283660 3788 283666 3800
rect 285398 3788 285404 3800
rect 283660 3760 285404 3788
rect 283660 3748 283666 3760
rect 285398 3748 285404 3760
rect 285456 3748 285462 3800
rect 287098 3748 287104 3800
rect 287156 3788 287162 3800
rect 288986 3788 288992 3800
rect 287156 3760 288992 3788
rect 287156 3748 287162 3760
rect 288986 3748 288992 3760
rect 289044 3748 289050 3800
rect 291698 3748 291704 3800
rect 291756 3788 291762 3800
rect 293678 3788 293684 3800
rect 291756 3760 293684 3788
rect 291756 3748 291762 3760
rect 293678 3748 293684 3760
rect 293736 3748 293742 3800
rect 294090 3748 294096 3800
rect 294148 3788 294154 3800
rect 296070 3788 296076 3800
rect 294148 3760 296076 3788
rect 294148 3748 294154 3760
rect 296070 3748 296076 3760
rect 296128 3748 296134 3800
rect 298690 3748 298696 3800
rect 298748 3788 298754 3800
rect 300762 3788 300768 3800
rect 298748 3760 300768 3788
rect 298748 3748 298754 3760
rect 300762 3748 300768 3760
rect 300820 3748 300826 3800
rect 300990 3748 300996 3800
rect 301048 3788 301054 3800
rect 303154 3788 303160 3800
rect 301048 3760 303160 3788
rect 301048 3748 301054 3760
rect 303154 3748 303160 3760
rect 303212 3748 303218 3800
rect 307982 3748 307988 3800
rect 308040 3788 308046 3800
rect 310238 3788 310244 3800
rect 308040 3760 310244 3788
rect 308040 3748 308046 3760
rect 310238 3748 310244 3760
rect 310296 3748 310302 3800
rect 316078 3748 316084 3800
rect 316136 3788 316142 3800
rect 318518 3788 318524 3800
rect 316136 3760 318524 3788
rect 316136 3748 316142 3760
rect 318518 3748 318524 3760
rect 318576 3748 318582 3800
rect 323070 3748 323076 3800
rect 323128 3788 323134 3800
rect 325602 3788 325608 3800
rect 323128 3760 325608 3788
rect 323128 3748 323134 3760
rect 325602 3748 325608 3760
rect 325660 3748 325666 3800
rect 63218 3000 63224 3052
rect 63276 3040 63282 3052
rect 65518 3040 65524 3052
rect 63276 3012 65524 3040
rect 63276 3000 63282 3012
rect 65518 3000 65524 3012
rect 65576 3000 65582 3052
rect 4062 2864 4068 2916
rect 4120 2904 4126 2916
rect 7466 2904 7472 2916
rect 4120 2876 7472 2904
rect 4120 2864 4126 2876
rect 7466 2864 7472 2876
rect 7524 2864 7530 2916
rect 18230 2864 18236 2916
rect 18288 2904 18294 2916
rect 21450 2904 21456 2916
rect 18288 2876 21456 2904
rect 18288 2864 18294 2876
rect 21450 2864 21456 2876
rect 21508 2864 21514 2916
rect 253382 2864 253388 2916
rect 253440 2904 253446 2916
rect 254670 2904 254676 2916
rect 253440 2876 254676 2904
rect 253440 2864 253446 2876
rect 254670 2864 254676 2876
rect 254728 2864 254734 2916
rect 6454 2796 6460 2848
rect 6512 2836 6518 2848
rect 9858 2836 9864 2848
rect 6512 2808 9864 2836
rect 6512 2796 6518 2808
rect 9858 2796 9864 2808
rect 9916 2796 9922 2848
rect 9950 2796 9956 2848
rect 10008 2836 10014 2848
rect 13262 2836 13268 2848
rect 10008 2808 13268 2836
rect 10008 2796 10014 2808
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 17034 2796 17040 2848
rect 17092 2836 17098 2848
rect 20254 2836 20260 2848
rect 17092 2808 20260 2836
rect 17092 2796 17098 2808
rect 20254 2796 20260 2808
rect 20312 2796 20318 2848
rect 28902 2796 28908 2848
rect 28960 2836 28966 2848
rect 31846 2836 31852 2848
rect 28960 2808 31852 2836
rect 28960 2796 28966 2808
rect 31846 2796 31852 2808
rect 31904 2796 31910 2848
rect 35986 2796 35992 2848
rect 36044 2836 36050 2848
rect 38838 2836 38844 2848
rect 36044 2808 38844 2836
rect 36044 2796 36050 2808
rect 38838 2796 38844 2808
rect 38896 2796 38902 2848
rect 39574 2796 39580 2848
rect 39632 2836 39638 2848
rect 42334 2836 42340 2848
rect 39632 2808 42340 2836
rect 39632 2796 39638 2808
rect 42334 2796 42340 2808
rect 42392 2796 42398 2848
rect 62022 2796 62028 2848
rect 62080 2836 62086 2848
rect 64414 2836 64420 2848
rect 62080 2808 64420 2836
rect 62080 2796 62086 2808
rect 64414 2796 64420 2808
rect 64472 2796 64478 2848
rect 65518 2796 65524 2848
rect 65576 2836 65582 2848
rect 67818 2836 67824 2848
rect 65576 2808 67824 2836
rect 65576 2796 65582 2808
rect 67818 2796 67824 2808
rect 67876 2796 67882 2848
rect 248874 2796 248880 2848
rect 248932 2836 248938 2848
rect 249978 2836 249984 2848
rect 248932 2808 249984 2836
rect 248932 2796 248938 2808
rect 249978 2796 249984 2808
rect 250036 2796 250042 2848
rect 251082 2796 251088 2848
rect 251140 2836 251146 2848
rect 252370 2836 252376 2848
rect 251140 2808 252376 2836
rect 251140 2796 251146 2808
rect 252370 2796 252376 2808
rect 252428 2796 252434 2848
rect 254578 2796 254584 2848
rect 254636 2836 254642 2848
rect 255866 2836 255872 2848
rect 254636 2808 255872 2836
rect 254636 2796 254642 2808
rect 255866 2796 255872 2808
rect 255924 2796 255930 2848
rect 309226 2796 309232 2848
rect 309284 2836 309290 2848
rect 311434 2836 311440 2848
rect 309284 2808 311440 2836
rect 309284 2796 309290 2808
rect 311434 2796 311440 2808
rect 311492 2796 311498 2848
rect 315022 2796 315028 2848
rect 315080 2836 315086 2848
rect 317322 2836 317328 2848
rect 315080 2808 317328 2836
rect 315080 2796 315086 2808
rect 317322 2796 317328 2808
rect 317380 2796 317386 2848
rect 411162 2796 411168 2848
rect 411220 2836 411226 2848
rect 415486 2836 415492 2848
rect 411220 2808 415492 2836
rect 411220 2796 411226 2808
rect 415486 2796 415492 2808
rect 415544 2796 415550 2848
rect 440142 2796 440148 2848
rect 440200 2836 440206 2848
rect 445018 2836 445024 2848
rect 440200 2808 445024 2836
rect 440200 2796 440206 2808
rect 445018 2796 445024 2808
rect 445076 2796 445082 2848
rect 449526 2796 449532 2848
rect 449584 2836 449590 2848
rect 454494 2836 454500 2848
rect 449584 2808 454500 2836
rect 449584 2796 449590 2808
rect 454494 2796 454500 2808
rect 454552 2796 454558 2848
rect 478506 2796 478512 2848
rect 478564 2836 478570 2848
rect 484026 2836 484032 2848
rect 478564 2808 484032 2836
rect 478564 2796 478570 2808
rect 484026 2796 484032 2808
rect 484084 2796 484090 2848
rect 487798 2796 487804 2848
rect 487856 2836 487862 2848
rect 493502 2836 493508 2848
rect 487856 2808 493508 2836
rect 487856 2796 487862 2808
rect 493502 2796 493508 2808
rect 493560 2796 493566 2848
rect 3234 1300 3240 1352
rect 3292 1340 3298 1352
rect 6362 1340 6368 1352
rect 3292 1312 6368 1340
rect 3292 1300 3298 1312
rect 6362 1300 6368 1312
rect 6420 1300 6426 1352
rect 60826 1300 60832 1352
rect 60884 1340 60890 1352
rect 63310 1340 63316 1352
rect 60884 1312 63316 1340
rect 60884 1300 60890 1312
rect 63310 1300 63316 1312
rect 63368 1300 63374 1352
rect 67910 1300 67916 1352
rect 67968 1340 67974 1352
rect 70118 1340 70124 1352
rect 67968 1312 70124 1340
rect 67968 1300 67974 1312
rect 70118 1300 70124 1312
rect 70176 1300 70182 1352
rect 76190 1300 76196 1352
rect 76248 1340 76254 1352
rect 78214 1340 78220 1352
rect 76248 1312 78220 1340
rect 76248 1300 76254 1312
rect 78214 1300 78220 1312
rect 78272 1300 78278 1352
rect 83274 1300 83280 1352
rect 83332 1340 83338 1352
rect 85206 1340 85212 1352
rect 83332 1312 85212 1340
rect 83332 1300 83338 1312
rect 85206 1300 85212 1312
rect 85264 1300 85270 1352
rect 85666 1300 85672 1352
rect 85724 1340 85730 1352
rect 87506 1340 87512 1352
rect 85724 1312 87512 1340
rect 85724 1300 85730 1312
rect 87506 1300 87512 1312
rect 87564 1300 87570 1352
rect 89162 1300 89168 1352
rect 89220 1340 89226 1352
rect 91002 1340 91008 1352
rect 89220 1312 91008 1340
rect 89220 1300 89226 1312
rect 91002 1300 91008 1312
rect 91060 1300 91066 1352
rect 91554 1300 91560 1352
rect 91612 1340 91618 1352
rect 93302 1340 93308 1352
rect 91612 1312 93308 1340
rect 91612 1300 91618 1312
rect 93302 1300 93308 1312
rect 93360 1300 93366 1352
rect 93946 1300 93952 1352
rect 94004 1340 94010 1352
rect 95694 1340 95700 1352
rect 94004 1312 95700 1340
rect 94004 1300 94010 1312
rect 95694 1300 95700 1312
rect 95752 1300 95758 1352
rect 97442 1300 97448 1352
rect 97500 1340 97506 1352
rect 99098 1340 99104 1352
rect 97500 1312 99104 1340
rect 97500 1300 97506 1312
rect 99098 1300 99104 1312
rect 99156 1300 99162 1352
rect 101030 1300 101036 1352
rect 101088 1340 101094 1352
rect 102594 1340 102600 1352
rect 101088 1312 102600 1340
rect 101088 1300 101094 1312
rect 102594 1300 102600 1312
rect 102652 1300 102658 1352
rect 104526 1300 104532 1352
rect 104584 1340 104590 1352
rect 106090 1340 106096 1352
rect 104584 1312 106096 1340
rect 104584 1300 104590 1312
rect 106090 1300 106096 1312
rect 106148 1300 106154 1352
rect 106918 1300 106924 1352
rect 106976 1340 106982 1352
rect 108390 1340 108396 1352
rect 106976 1312 108396 1340
rect 106976 1300 106982 1312
rect 108390 1300 108396 1312
rect 108448 1300 108454 1352
rect 109310 1300 109316 1352
rect 109368 1340 109374 1352
rect 110690 1340 110696 1352
rect 109368 1312 110696 1340
rect 109368 1300 109374 1312
rect 110690 1300 110696 1312
rect 110748 1300 110754 1352
rect 112806 1300 112812 1352
rect 112864 1340 112870 1352
rect 114186 1340 114192 1352
rect 112864 1312 114192 1340
rect 112864 1300 112870 1312
rect 114186 1300 114192 1312
rect 114244 1300 114250 1352
rect 116394 1300 116400 1352
rect 116452 1340 116458 1352
rect 117682 1340 117688 1352
rect 116452 1312 117688 1340
rect 116452 1300 116458 1312
rect 117682 1300 117688 1312
rect 117740 1300 117746 1352
rect 119890 1300 119896 1352
rect 119948 1340 119954 1352
rect 121178 1340 121184 1352
rect 119948 1312 121184 1340
rect 119948 1300 119954 1312
rect 121178 1300 121184 1312
rect 121236 1300 121242 1352
rect 125870 1300 125876 1352
rect 125928 1340 125934 1352
rect 126974 1340 126980 1352
rect 125928 1312 126980 1340
rect 125928 1300 125934 1312
rect 126974 1300 126980 1312
rect 127032 1300 127038 1352
rect 129366 1300 129372 1352
rect 129424 1340 129430 1352
rect 130470 1340 130476 1352
rect 129424 1312 130476 1340
rect 129424 1300 129430 1312
rect 130470 1300 130476 1312
rect 130528 1300 130534 1352
rect 130562 1300 130568 1352
rect 130620 1340 130626 1352
rect 131574 1340 131580 1352
rect 130620 1312 131580 1340
rect 130620 1300 130626 1312
rect 131574 1300 131580 1312
rect 131632 1300 131638 1352
rect 131758 1300 131764 1352
rect 131816 1340 131822 1352
rect 132770 1340 132776 1352
rect 131816 1312 132776 1340
rect 131816 1300 131822 1312
rect 132770 1300 132776 1312
rect 132828 1300 132834 1352
rect 132954 1300 132960 1352
rect 133012 1340 133018 1352
rect 133966 1340 133972 1352
rect 133012 1312 133972 1340
rect 133012 1300 133018 1312
rect 133966 1300 133972 1312
rect 134024 1300 134030 1352
rect 137646 1300 137652 1352
rect 137704 1340 137710 1352
rect 138566 1340 138572 1352
rect 137704 1312 138572 1340
rect 137704 1300 137710 1312
rect 138566 1300 138572 1312
rect 138624 1300 138630 1352
rect 144730 1300 144736 1352
rect 144788 1340 144794 1352
rect 145558 1340 145564 1352
rect 144788 1312 145564 1340
rect 144788 1300 144794 1312
rect 145558 1300 145564 1312
rect 145616 1300 145622 1352
rect 145926 1300 145932 1352
rect 145984 1340 145990 1352
rect 146662 1340 146668 1352
rect 145984 1312 146668 1340
rect 145984 1300 145990 1312
rect 146662 1300 146668 1312
rect 146720 1300 146726 1352
rect 148318 1300 148324 1352
rect 148376 1340 148382 1352
rect 149054 1340 149060 1352
rect 148376 1312 149060 1340
rect 148376 1300 148382 1312
rect 149054 1300 149060 1312
rect 149112 1300 149118 1352
rect 154206 1300 154212 1352
rect 154264 1340 154270 1352
rect 154850 1340 154856 1352
rect 154264 1312 154856 1340
rect 154264 1300 154270 1312
rect 154850 1300 154856 1312
rect 154908 1300 154914 1352
rect 162486 1300 162492 1352
rect 162544 1340 162550 1352
rect 162946 1340 162952 1352
rect 162544 1312 162952 1340
rect 162544 1300 162550 1312
rect 162946 1300 162952 1312
rect 163004 1300 163010 1352
rect 266262 1300 266268 1352
rect 266320 1340 266326 1352
rect 267734 1340 267740 1352
rect 266320 1312 267740 1340
rect 266320 1300 266326 1312
rect 267734 1300 267740 1312
rect 267792 1300 267798 1352
rect 273162 1300 273168 1352
rect 273220 1340 273226 1352
rect 274818 1340 274824 1352
rect 273220 1312 274824 1340
rect 273220 1300 273226 1312
rect 274818 1300 274824 1312
rect 274876 1300 274882 1352
rect 280062 1300 280068 1352
rect 280120 1340 280126 1352
rect 281902 1340 281908 1352
rect 280120 1312 281908 1340
rect 280120 1300 280126 1312
rect 281902 1300 281908 1312
rect 281960 1300 281966 1352
rect 282546 1300 282552 1352
rect 282604 1340 282610 1352
rect 284294 1340 284300 1352
rect 282604 1312 284300 1340
rect 282604 1300 282610 1312
rect 284294 1300 284300 1312
rect 284352 1300 284358 1352
rect 288342 1300 288348 1352
rect 288400 1340 288406 1352
rect 290182 1340 290188 1352
rect 288400 1312 290188 1340
rect 288400 1300 288406 1312
rect 290182 1300 290188 1312
rect 290240 1300 290246 1352
rect 295242 1300 295248 1352
rect 295300 1340 295306 1352
rect 297266 1340 297272 1352
rect 295300 1312 297272 1340
rect 295300 1300 295306 1312
rect 297266 1300 297272 1312
rect 297324 1300 297330 1352
rect 297542 1300 297548 1352
rect 297600 1340 297606 1352
rect 299658 1340 299664 1352
rect 297600 1312 299664 1340
rect 297600 1300 297606 1312
rect 299658 1300 299664 1312
rect 299716 1300 299722 1352
rect 302142 1300 302148 1352
rect 302200 1340 302206 1352
rect 304350 1340 304356 1352
rect 302200 1312 304356 1340
rect 302200 1300 302206 1312
rect 304350 1300 304356 1312
rect 304408 1300 304414 1352
rect 305730 1300 305736 1352
rect 305788 1340 305794 1352
rect 307938 1340 307944 1352
rect 305788 1312 307944 1340
rect 305788 1300 305794 1312
rect 307938 1300 307944 1312
rect 307996 1300 308002 1352
rect 310330 1300 310336 1352
rect 310388 1340 310394 1352
rect 312630 1340 312636 1352
rect 310388 1312 312636 1340
rect 310388 1300 310394 1312
rect 312630 1300 312636 1312
rect 312688 1300 312694 1352
rect 313826 1300 313832 1352
rect 313884 1340 313890 1352
rect 316218 1340 316224 1352
rect 313884 1312 316224 1340
rect 313884 1300 313890 1312
rect 316218 1300 316224 1312
rect 316276 1300 316282 1352
rect 317230 1300 317236 1352
rect 317288 1340 317294 1352
rect 319714 1340 319720 1352
rect 317288 1312 319720 1340
rect 317288 1300 317294 1312
rect 319714 1300 319720 1312
rect 319772 1300 319778 1352
rect 321922 1300 321928 1352
rect 321980 1340 321986 1352
rect 324406 1340 324412 1352
rect 321980 1312 324412 1340
rect 321980 1300 321986 1312
rect 324406 1300 324412 1312
rect 324464 1300 324470 1352
rect 326614 1300 326620 1352
rect 326672 1340 326678 1352
rect 329190 1340 329196 1352
rect 326672 1312 329196 1340
rect 326672 1300 326678 1312
rect 329190 1300 329196 1312
rect 329248 1300 329254 1352
rect 332410 1300 332416 1352
rect 332468 1340 332474 1352
rect 335078 1340 335084 1352
rect 332468 1312 335084 1340
rect 332468 1300 332474 1312
rect 335078 1300 335084 1312
rect 335136 1300 335142 1352
rect 335906 1300 335912 1352
rect 335964 1340 335970 1352
rect 338666 1340 338672 1352
rect 335964 1312 338672 1340
rect 335964 1300 335970 1312
rect 338666 1300 338672 1312
rect 338724 1300 338730 1352
rect 339310 1300 339316 1352
rect 339368 1340 339374 1352
rect 342162 1340 342168 1352
rect 339368 1312 342168 1340
rect 339368 1300 339374 1312
rect 342162 1300 342168 1312
rect 342220 1300 342226 1352
rect 345106 1300 345112 1352
rect 345164 1340 345170 1352
rect 348050 1340 348056 1352
rect 345164 1312 348056 1340
rect 345164 1300 345170 1312
rect 348050 1300 348056 1312
rect 348108 1300 348114 1352
rect 349798 1300 349804 1352
rect 349856 1340 349862 1352
rect 352834 1340 352840 1352
rect 349856 1312 352840 1340
rect 349856 1300 349862 1312
rect 352834 1300 352840 1312
rect 352892 1300 352898 1352
rect 353202 1300 353208 1352
rect 353260 1340 353266 1352
rect 356330 1340 356336 1352
rect 353260 1312 356336 1340
rect 353260 1300 353266 1312
rect 356330 1300 356336 1312
rect 356388 1300 356394 1352
rect 356698 1300 356704 1352
rect 356756 1340 356762 1352
rect 359918 1340 359924 1352
rect 356756 1312 359924 1340
rect 356756 1300 356762 1312
rect 359918 1300 359924 1312
rect 359976 1300 359982 1352
rect 362586 1300 362592 1352
rect 362644 1340 362650 1352
rect 365806 1340 365812 1352
rect 362644 1312 365812 1340
rect 362644 1300 362650 1312
rect 365806 1300 365812 1312
rect 365864 1300 365870 1352
rect 367186 1300 367192 1352
rect 367244 1340 367250 1352
rect 370590 1340 370596 1352
rect 367244 1312 370596 1340
rect 367244 1300 367250 1312
rect 370590 1300 370596 1312
rect 370648 1300 370654 1352
rect 370682 1300 370688 1352
rect 370740 1340 370746 1352
rect 374086 1340 374092 1352
rect 370740 1312 374092 1340
rect 370740 1300 370746 1312
rect 374086 1300 374092 1312
rect 374144 1300 374150 1352
rect 376386 1300 376392 1352
rect 376444 1340 376450 1352
rect 379974 1340 379980 1352
rect 376444 1312 379980 1340
rect 376444 1300 376450 1312
rect 379974 1300 379980 1312
rect 380032 1300 380038 1352
rect 385770 1300 385776 1352
rect 385828 1340 385834 1352
rect 389450 1340 389456 1352
rect 385828 1312 389456 1340
rect 385828 1300 385834 1312
rect 389450 1300 389456 1312
rect 389508 1300 389514 1352
rect 395062 1300 395068 1352
rect 395120 1340 395126 1352
rect 398926 1340 398932 1352
rect 395120 1312 398932 1340
rect 395120 1300 395126 1312
rect 398926 1300 398932 1312
rect 398984 1300 398990 1352
rect 399662 1300 399668 1352
rect 399720 1340 399726 1352
rect 403618 1340 403624 1352
rect 399720 1312 403624 1340
rect 399720 1300 399726 1312
rect 403618 1300 403624 1312
rect 403676 1300 403682 1352
rect 405458 1300 405464 1352
rect 405516 1340 405522 1352
rect 409598 1340 409604 1352
rect 405516 1312 409604 1340
rect 405516 1300 405522 1312
rect 409598 1300 409604 1312
rect 409656 1300 409662 1352
rect 413554 1300 413560 1352
rect 413612 1340 413618 1352
rect 417878 1340 417884 1352
rect 413612 1312 417884 1340
rect 413612 1300 413618 1312
rect 417878 1300 417884 1312
rect 417936 1300 417942 1352
rect 422846 1300 422852 1352
rect 422904 1340 422910 1352
rect 427262 1340 427268 1352
rect 422904 1312 427268 1340
rect 422904 1300 422910 1312
rect 427262 1300 427268 1312
rect 427320 1300 427326 1352
rect 427538 1300 427544 1352
rect 427596 1340 427602 1352
rect 431862 1340 431868 1352
rect 427596 1312 431868 1340
rect 427596 1300 427602 1312
rect 431862 1300 431868 1312
rect 431920 1300 431926 1352
rect 433242 1300 433248 1352
rect 433300 1340 433306 1352
rect 437842 1340 437848 1352
rect 433300 1312 437848 1340
rect 433300 1300 433306 1312
rect 437842 1300 437848 1312
rect 437900 1300 437906 1352
rect 441430 1300 441436 1352
rect 441488 1340 441494 1352
rect 445846 1340 445852 1352
rect 441488 1312 445852 1340
rect 441488 1300 441494 1312
rect 445846 1300 445852 1312
rect 445904 1300 445910 1352
rect 447226 1300 447232 1352
rect 447284 1340 447290 1352
rect 452102 1340 452108 1352
rect 447284 1312 452108 1340
rect 447284 1300 447290 1312
rect 452102 1300 452108 1312
rect 452160 1300 452166 1352
rect 453022 1300 453028 1352
rect 453080 1340 453086 1352
rect 458082 1340 458088 1352
rect 453080 1312 458088 1340
rect 453080 1300 453086 1312
rect 458082 1300 458088 1312
rect 458140 1300 458146 1352
rect 458818 1300 458824 1352
rect 458876 1340 458882 1352
rect 463970 1340 463976 1352
rect 458876 1312 463976 1340
rect 458876 1300 458882 1312
rect 463970 1300 463976 1312
rect 464028 1300 464034 1352
rect 471606 1300 471612 1352
rect 471664 1340 471670 1352
rect 476574 1340 476580 1352
rect 471664 1312 476580 1340
rect 471664 1300 471670 1312
rect 476574 1300 476580 1312
rect 476632 1300 476638 1352
rect 477402 1300 477408 1352
rect 477460 1340 477466 1352
rect 482462 1340 482468 1352
rect 477460 1312 482468 1340
rect 477460 1300 477466 1312
rect 482462 1300 482468 1312
rect 482520 1300 482526 1352
rect 483198 1300 483204 1352
rect 483256 1340 483262 1352
rect 488810 1340 488816 1352
rect 483256 1312 488816 1340
rect 483256 1300 483262 1312
rect 488810 1300 488816 1312
rect 488868 1300 488874 1352
rect 490098 1300 490104 1352
rect 490156 1340 490162 1352
rect 495526 1340 495532 1352
rect 490156 1312 495532 1340
rect 490156 1300 490162 1312
rect 495526 1300 495532 1312
rect 495584 1300 495590 1352
rect 497090 1300 497096 1352
rect 497148 1340 497154 1352
rect 502978 1340 502984 1352
rect 497148 1312 502984 1340
rect 497148 1300 497154 1312
rect 502978 1300 502984 1312
rect 503036 1300 503042 1352
rect 504082 1300 504088 1352
rect 504140 1340 504146 1352
rect 509694 1340 509700 1352
rect 504140 1312 509700 1340
rect 504140 1300 504146 1312
rect 509694 1300 509700 1312
rect 509752 1300 509758 1352
rect 509878 1300 509884 1352
rect 509936 1340 509942 1352
rect 515766 1340 515772 1352
rect 509936 1312 515772 1340
rect 509936 1300 509942 1312
rect 515766 1300 515772 1312
rect 515824 1300 515830 1352
rect 519170 1300 519176 1352
rect 519228 1340 519234 1352
rect 525426 1340 525432 1352
rect 519228 1312 525432 1340
rect 519228 1300 519234 1312
rect 525426 1300 525432 1312
rect 525484 1300 525490 1352
rect 526070 1300 526076 1352
rect 526128 1340 526134 1352
rect 532142 1340 532148 1352
rect 526128 1312 532148 1340
rect 526128 1300 526134 1312
rect 532142 1300 532148 1312
rect 532200 1300 532206 1352
rect 534258 1300 534264 1352
rect 534316 1340 534322 1352
rect 540422 1340 540428 1352
rect 534316 1312 540428 1340
rect 534316 1300 534322 1312
rect 540422 1300 540428 1312
rect 540480 1300 540486 1352
rect 542262 1300 542268 1352
rect 542320 1340 542326 1352
rect 549070 1340 549076 1352
rect 542320 1312 549076 1340
rect 542320 1300 542326 1312
rect 549070 1300 549076 1312
rect 549128 1300 549134 1352
rect 551646 1300 551652 1352
rect 551704 1340 551710 1352
rect 558546 1340 558552 1352
rect 551704 1312 558552 1340
rect 551704 1300 551710 1312
rect 558546 1300 558552 1312
rect 558604 1300 558610 1352
rect 560938 1300 560944 1352
rect 560996 1340 561002 1352
rect 568022 1340 568028 1352
rect 560996 1312 568028 1340
rect 560996 1300 561002 1312
rect 568022 1300 568028 1312
rect 568080 1300 568086 1352
rect 571242 1300 571248 1352
rect 571300 1340 571306 1352
rect 578602 1340 578608 1352
rect 571300 1312 578608 1340
rect 571300 1300 571306 1312
rect 578602 1300 578608 1312
rect 578660 1300 578666 1352
rect 74994 1232 75000 1284
rect 75052 1272 75058 1284
rect 77110 1272 77116 1284
rect 75052 1244 77116 1272
rect 75052 1232 75058 1244
rect 77110 1232 77116 1244
rect 77168 1232 77174 1284
rect 77386 1232 77392 1284
rect 77444 1272 77450 1284
rect 79410 1272 79416 1284
rect 77444 1244 79416 1272
rect 77444 1232 77450 1244
rect 79410 1232 79416 1244
rect 79468 1232 79474 1284
rect 82078 1232 82084 1284
rect 82136 1272 82142 1284
rect 84010 1272 84016 1284
rect 82136 1244 84016 1272
rect 82136 1232 82142 1244
rect 84010 1232 84016 1244
rect 84068 1232 84074 1284
rect 84470 1232 84476 1284
rect 84528 1272 84534 1284
rect 86402 1272 86408 1284
rect 84528 1244 86408 1272
rect 84528 1232 84534 1244
rect 86402 1232 86408 1244
rect 86460 1232 86466 1284
rect 90358 1232 90364 1284
rect 90416 1272 90422 1284
rect 92198 1272 92204 1284
rect 90416 1244 92204 1272
rect 90416 1232 90422 1244
rect 92198 1232 92204 1244
rect 92256 1232 92262 1284
rect 92750 1232 92756 1284
rect 92808 1272 92814 1284
rect 94498 1272 94504 1284
rect 92808 1244 94504 1272
rect 92808 1232 92814 1244
rect 94498 1232 94504 1244
rect 94556 1232 94562 1284
rect 98638 1232 98644 1284
rect 98696 1272 98702 1284
rect 100294 1272 100300 1284
rect 98696 1244 100300 1272
rect 98696 1232 98702 1244
rect 100294 1232 100300 1244
rect 100352 1232 100358 1284
rect 102226 1232 102232 1284
rect 102284 1272 102290 1284
rect 103790 1272 103796 1284
rect 102284 1244 103796 1272
rect 102284 1232 102290 1244
rect 103790 1232 103796 1244
rect 103848 1232 103854 1284
rect 108114 1232 108120 1284
rect 108172 1272 108178 1284
rect 109586 1272 109592 1284
rect 108172 1244 109592 1272
rect 108172 1232 108178 1244
rect 109586 1232 109592 1244
rect 109644 1232 109650 1284
rect 110506 1232 110512 1284
rect 110564 1272 110570 1284
rect 111886 1272 111892 1284
rect 110564 1244 111892 1272
rect 110564 1232 110570 1244
rect 111886 1232 111892 1244
rect 111944 1232 111950 1284
rect 115198 1232 115204 1284
rect 115256 1272 115262 1284
rect 116578 1272 116584 1284
rect 115256 1244 116584 1272
rect 115256 1232 115262 1244
rect 116578 1232 116584 1244
rect 116636 1232 116642 1284
rect 117590 1232 117596 1284
rect 117648 1272 117654 1284
rect 118878 1272 118884 1284
rect 117648 1244 118884 1272
rect 117648 1232 117654 1244
rect 118878 1232 118884 1244
rect 118936 1232 118942 1284
rect 122282 1232 122288 1284
rect 122340 1272 122346 1284
rect 123478 1272 123484 1284
rect 122340 1244 123484 1272
rect 122340 1232 122346 1244
rect 123478 1232 123484 1244
rect 123536 1232 123542 1284
rect 124674 1232 124680 1284
rect 124732 1272 124738 1284
rect 125778 1272 125784 1284
rect 124732 1244 125784 1272
rect 124732 1232 124738 1244
rect 125778 1232 125784 1244
rect 125836 1232 125842 1284
rect 128170 1232 128176 1284
rect 128228 1272 128234 1284
rect 129274 1272 129280 1284
rect 128228 1244 129280 1272
rect 128228 1232 128234 1244
rect 129274 1232 129280 1244
rect 129332 1232 129338 1284
rect 136450 1232 136456 1284
rect 136508 1272 136514 1284
rect 137370 1272 137376 1284
rect 136508 1244 137376 1272
rect 136508 1232 136514 1244
rect 137370 1232 137376 1244
rect 137428 1232 137434 1284
rect 138842 1232 138848 1284
rect 138900 1272 138906 1284
rect 139762 1272 139768 1284
rect 138900 1244 139768 1272
rect 138900 1232 138906 1244
rect 139762 1232 139768 1244
rect 139820 1232 139826 1284
rect 140038 1232 140044 1284
rect 140096 1272 140102 1284
rect 140866 1272 140872 1284
rect 140096 1244 140872 1272
rect 140096 1232 140102 1244
rect 140866 1232 140872 1244
rect 140924 1232 140930 1284
rect 281350 1232 281356 1284
rect 281408 1272 281414 1284
rect 283098 1272 283104 1284
rect 281408 1244 283104 1272
rect 281408 1232 281414 1244
rect 283098 1232 283104 1244
rect 283156 1232 283162 1284
rect 289446 1232 289452 1284
rect 289504 1272 289510 1284
rect 291378 1272 291384 1284
rect 289504 1244 291384 1272
rect 289504 1232 289510 1244
rect 291378 1232 291384 1244
rect 291436 1232 291442 1284
rect 296438 1232 296444 1284
rect 296496 1272 296502 1284
rect 298462 1272 298468 1284
rect 296496 1244 298468 1272
rect 296496 1232 296502 1244
rect 298462 1232 298468 1244
rect 298520 1232 298526 1284
rect 303338 1232 303344 1284
rect 303396 1272 303402 1284
rect 305546 1272 305552 1284
rect 303396 1244 305552 1272
rect 303396 1232 303402 1244
rect 305546 1232 305552 1244
rect 305604 1232 305610 1284
rect 312538 1232 312544 1284
rect 312596 1272 312602 1284
rect 315022 1272 315028 1284
rect 312596 1244 315028 1272
rect 312596 1232 312602 1244
rect 315022 1232 315028 1244
rect 315080 1232 315086 1284
rect 318426 1232 318432 1284
rect 318484 1272 318490 1284
rect 320910 1272 320916 1284
rect 318484 1244 320916 1272
rect 318484 1232 318490 1244
rect 320910 1232 320916 1244
rect 320968 1232 320974 1284
rect 328914 1232 328920 1284
rect 328972 1272 328978 1284
rect 331582 1272 331588 1284
rect 328972 1244 331588 1272
rect 328972 1232 328978 1244
rect 331582 1232 331588 1244
rect 331640 1232 331646 1284
rect 334710 1232 334716 1284
rect 334768 1272 334774 1284
rect 337470 1272 337476 1284
rect 334768 1244 337476 1272
rect 334768 1232 334774 1244
rect 337470 1232 337476 1244
rect 337528 1232 337534 1284
rect 340506 1232 340512 1284
rect 340564 1272 340570 1284
rect 343358 1272 343364 1284
rect 340564 1244 343364 1272
rect 340564 1232 340570 1244
rect 343358 1232 343364 1244
rect 343416 1232 343422 1284
rect 344002 1232 344008 1284
rect 344060 1272 344066 1284
rect 346946 1272 346952 1284
rect 344060 1244 346952 1272
rect 344060 1232 344066 1244
rect 346946 1232 346952 1244
rect 347004 1232 347010 1284
rect 348602 1232 348608 1284
rect 348660 1272 348666 1284
rect 351638 1272 351644 1284
rect 348660 1244 351644 1272
rect 348660 1232 348666 1244
rect 351638 1232 351644 1244
rect 351696 1232 351702 1284
rect 352098 1232 352104 1284
rect 352156 1272 352162 1284
rect 355226 1272 355232 1284
rect 352156 1244 355232 1272
rect 352156 1232 352162 1244
rect 355226 1232 355232 1244
rect 355284 1232 355290 1284
rect 355594 1232 355600 1284
rect 355652 1272 355658 1284
rect 358722 1272 358728 1284
rect 355652 1244 358728 1272
rect 355652 1232 355658 1244
rect 358722 1232 358728 1244
rect 358780 1232 358786 1284
rect 359090 1232 359096 1284
rect 359148 1272 359154 1284
rect 362310 1272 362316 1284
rect 359148 1244 362316 1272
rect 359148 1232 359154 1244
rect 362310 1232 362316 1244
rect 362368 1232 362374 1284
rect 363690 1232 363696 1284
rect 363748 1272 363754 1284
rect 367002 1272 367008 1284
rect 363748 1244 367008 1272
rect 363748 1232 363754 1244
rect 367002 1232 367008 1244
rect 367060 1232 367066 1284
rect 372982 1232 372988 1284
rect 373040 1272 373046 1284
rect 376478 1272 376484 1284
rect 373040 1244 376484 1272
rect 373040 1232 373046 1244
rect 376478 1232 376484 1244
rect 376536 1232 376542 1284
rect 377582 1232 377588 1284
rect 377640 1272 377646 1284
rect 381170 1272 381176 1284
rect 377640 1244 381176 1272
rect 377640 1232 377646 1244
rect 381170 1232 381176 1244
rect 381228 1232 381234 1284
rect 388070 1232 388076 1284
rect 388128 1272 388134 1284
rect 391842 1272 391848 1284
rect 388128 1244 391848 1272
rect 388128 1232 388134 1244
rect 391842 1232 391848 1244
rect 391900 1232 391906 1284
rect 393866 1232 393872 1284
rect 393924 1272 393930 1284
rect 397730 1272 397736 1284
rect 393924 1244 397736 1272
rect 393924 1232 393930 1244
rect 397730 1232 397736 1244
rect 397788 1232 397794 1284
rect 403158 1232 403164 1284
rect 403216 1272 403222 1284
rect 407206 1272 407212 1284
rect 403216 1244 407212 1272
rect 403216 1232 403222 1244
rect 407206 1232 407212 1244
rect 407264 1232 407270 1284
rect 410058 1232 410064 1284
rect 410116 1272 410122 1284
rect 414290 1272 414296 1284
rect 410116 1244 414296 1272
rect 410116 1232 410122 1244
rect 414290 1232 414296 1244
rect 414348 1232 414354 1284
rect 418246 1232 418252 1284
rect 418304 1272 418310 1284
rect 422570 1272 422576 1284
rect 418304 1244 422576 1272
rect 418304 1232 418310 1244
rect 422570 1232 422576 1244
rect 422628 1232 422634 1284
rect 426342 1232 426348 1284
rect 426400 1272 426406 1284
rect 430850 1272 430856 1284
rect 426400 1244 430856 1272
rect 426400 1232 426406 1244
rect 430850 1232 430856 1244
rect 430908 1232 430914 1284
rect 435634 1232 435640 1284
rect 435692 1272 435698 1284
rect 439958 1272 439964 1284
rect 435692 1244 439964 1272
rect 435692 1232 435698 1244
rect 439958 1232 439964 1244
rect 440016 1232 440022 1284
rect 442626 1232 442632 1284
rect 442684 1272 442690 1284
rect 447410 1272 447416 1284
rect 442684 1244 447416 1272
rect 442684 1232 442690 1244
rect 447410 1232 447416 1244
rect 447468 1232 447474 1284
rect 457622 1232 457628 1284
rect 457680 1272 457686 1284
rect 462406 1272 462412 1284
rect 457680 1244 462412 1272
rect 457680 1232 457686 1244
rect 462406 1232 462412 1244
rect 462464 1232 462470 1284
rect 468110 1232 468116 1284
rect 468168 1272 468174 1284
rect 473078 1272 473084 1284
rect 468168 1244 473084 1272
rect 468168 1232 468174 1244
rect 473078 1232 473084 1244
rect 473136 1232 473142 1284
rect 475102 1232 475108 1284
rect 475160 1272 475166 1284
rect 480530 1272 480536 1284
rect 475160 1244 480536 1272
rect 475160 1232 475166 1244
rect 480530 1232 480536 1244
rect 480588 1232 480594 1284
rect 485498 1232 485504 1284
rect 485556 1272 485562 1284
rect 490742 1272 490748 1284
rect 485556 1244 490748 1272
rect 485556 1232 485562 1244
rect 490742 1232 490748 1244
rect 490800 1232 490806 1284
rect 492490 1232 492496 1284
rect 492548 1272 492554 1284
rect 498194 1272 498200 1284
rect 492548 1244 498200 1272
rect 492548 1232 492554 1244
rect 498194 1232 498200 1244
rect 498252 1232 498258 1284
rect 498286 1232 498292 1284
rect 498344 1272 498350 1284
rect 503806 1272 503812 1284
rect 498344 1244 503812 1272
rect 498344 1232 498350 1244
rect 503806 1232 503812 1244
rect 503864 1232 503870 1284
rect 510982 1232 510988 1284
rect 511040 1272 511046 1284
rect 517146 1272 517152 1284
rect 511040 1244 517152 1272
rect 511040 1232 511046 1244
rect 517146 1232 517152 1244
rect 517204 1232 517210 1284
rect 517974 1232 517980 1284
rect 518032 1272 518038 1284
rect 523862 1272 523868 1284
rect 518032 1244 523868 1272
rect 518032 1232 518038 1244
rect 523862 1232 523868 1244
rect 523920 1232 523926 1284
rect 527266 1232 527272 1284
rect 527324 1272 527330 1284
rect 533706 1272 533712 1284
rect 527324 1244 533712 1272
rect 527324 1232 527330 1244
rect 533706 1232 533712 1244
rect 533764 1232 533770 1284
rect 541158 1232 541164 1284
rect 541216 1272 541222 1284
rect 547874 1272 547880 1284
rect 541216 1244 547880 1272
rect 541216 1232 541222 1244
rect 547874 1232 547880 1244
rect 547932 1232 547938 1284
rect 548150 1232 548156 1284
rect 548208 1272 548214 1284
rect 554958 1272 554964 1284
rect 548208 1244 554964 1272
rect 548208 1232 548214 1244
rect 554958 1232 554964 1244
rect 555016 1232 555022 1284
rect 562042 1232 562048 1284
rect 562100 1272 562106 1284
rect 569126 1272 569132 1284
rect 562100 1244 569132 1272
rect 562100 1232 562106 1244
rect 569126 1232 569132 1244
rect 569184 1232 569190 1284
rect 570138 1232 570144 1284
rect 570196 1272 570202 1284
rect 577406 1272 577412 1284
rect 570196 1244 577412 1272
rect 570196 1232 570202 1244
rect 577406 1232 577412 1244
rect 577464 1232 577470 1284
rect 99834 1164 99840 1216
rect 99892 1204 99898 1216
rect 101490 1204 101496 1216
rect 99892 1176 101496 1204
rect 99892 1164 99898 1176
rect 101490 1164 101496 1176
rect 101548 1164 101554 1216
rect 114002 1164 114008 1216
rect 114060 1204 114066 1216
rect 115382 1204 115388 1216
rect 114060 1176 115388 1204
rect 114060 1164 114066 1176
rect 115382 1164 115388 1176
rect 115440 1164 115446 1216
rect 311526 1164 311532 1216
rect 311584 1204 311590 1216
rect 313826 1204 313832 1216
rect 311584 1176 313832 1204
rect 311584 1164 311590 1176
rect 313826 1164 313832 1176
rect 313884 1164 313890 1216
rect 319622 1164 319628 1216
rect 319680 1204 319686 1216
rect 322106 1204 322112 1216
rect 319680 1176 322112 1204
rect 319680 1164 319686 1176
rect 322106 1164 322112 1176
rect 322164 1164 322170 1216
rect 330018 1164 330024 1216
rect 330076 1204 330082 1216
rect 332686 1204 332692 1216
rect 330076 1176 332692 1204
rect 330076 1164 330082 1176
rect 332686 1164 332692 1176
rect 332744 1164 332750 1216
rect 337010 1164 337016 1216
rect 337068 1204 337074 1216
rect 339862 1204 339868 1216
rect 337068 1176 339868 1204
rect 337068 1164 337074 1176
rect 339862 1164 339868 1176
rect 339920 1164 339926 1216
rect 341702 1164 341708 1216
rect 341760 1204 341766 1216
rect 344554 1204 344560 1216
rect 341760 1176 344560 1204
rect 341760 1164 341766 1176
rect 344554 1164 344560 1176
rect 344612 1164 344618 1216
rect 357894 1164 357900 1216
rect 357952 1204 357958 1216
rect 361114 1204 361120 1216
rect 357952 1176 361120 1204
rect 357952 1164 357958 1176
rect 361114 1164 361120 1176
rect 361172 1164 361178 1216
rect 364886 1164 364892 1216
rect 364944 1204 364950 1216
rect 368198 1204 368204 1216
rect 364944 1176 368204 1204
rect 364944 1164 364950 1176
rect 368198 1164 368204 1176
rect 368256 1164 368262 1216
rect 375282 1164 375288 1216
rect 375340 1204 375346 1216
rect 378870 1204 378876 1216
rect 375340 1176 378876 1204
rect 375340 1164 375346 1176
rect 378870 1164 378876 1176
rect 378928 1164 378934 1216
rect 381078 1164 381084 1216
rect 381136 1204 381142 1216
rect 384758 1204 384764 1216
rect 381136 1176 384764 1204
rect 381136 1164 381142 1176
rect 384758 1164 384764 1176
rect 384816 1164 384822 1216
rect 390370 1164 390376 1216
rect 390428 1204 390434 1216
rect 394234 1204 394240 1216
rect 390428 1176 394240 1204
rect 390428 1164 390434 1176
rect 394234 1164 394240 1176
rect 394292 1164 394298 1216
rect 396166 1164 396172 1216
rect 396224 1204 396230 1216
rect 400122 1204 400128 1216
rect 396224 1176 400128 1204
rect 396224 1164 396230 1176
rect 400122 1164 400128 1176
rect 400180 1164 400186 1216
rect 400858 1164 400864 1216
rect 400916 1204 400922 1216
rect 404814 1204 404820 1216
rect 400916 1176 404820 1204
rect 400916 1164 400922 1176
rect 404814 1164 404820 1176
rect 404872 1164 404878 1216
rect 407758 1164 407764 1216
rect 407816 1204 407822 1216
rect 411898 1204 411904 1216
rect 407816 1176 411904 1204
rect 407816 1164 407822 1176
rect 411898 1164 411904 1176
rect 411956 1164 411962 1216
rect 420546 1164 420552 1216
rect 420604 1204 420610 1216
rect 424962 1204 424968 1216
rect 420604 1176 424968 1204
rect 420604 1164 420610 1176
rect 424962 1164 424968 1176
rect 425020 1164 425026 1216
rect 425146 1164 425152 1216
rect 425204 1204 425210 1216
rect 429654 1204 429660 1216
rect 425204 1176 429660 1204
rect 425204 1164 425210 1176
rect 429654 1164 429660 1176
rect 429712 1164 429718 1216
rect 436738 1164 436744 1216
rect 436796 1204 436802 1216
rect 441522 1204 441528 1216
rect 436796 1176 441528 1204
rect 436796 1164 436802 1176
rect 441522 1164 441528 1176
rect 441580 1164 441586 1216
rect 444926 1164 444932 1216
rect 444984 1204 444990 1216
rect 449802 1204 449808 1216
rect 444984 1176 449808 1204
rect 444984 1164 444990 1176
rect 449802 1164 449808 1176
rect 449860 1164 449866 1216
rect 450722 1164 450728 1216
rect 450780 1204 450786 1216
rect 455690 1204 455696 1216
rect 450780 1176 455696 1204
rect 450780 1164 450786 1176
rect 455690 1164 455696 1176
rect 455748 1164 455754 1216
rect 456518 1164 456524 1216
rect 456576 1204 456582 1216
rect 461578 1204 461584 1216
rect 456576 1176 461584 1204
rect 456576 1164 456582 1176
rect 461578 1164 461584 1176
rect 461636 1164 461642 1216
rect 462222 1164 462228 1216
rect 462280 1204 462286 1216
rect 467466 1204 467472 1216
rect 462280 1176 467472 1204
rect 462280 1164 462286 1176
rect 467466 1164 467472 1176
rect 467524 1164 467530 1216
rect 472710 1164 472716 1216
rect 472768 1204 472774 1216
rect 478138 1204 478144 1216
rect 472768 1176 478144 1204
rect 472768 1164 472774 1176
rect 478138 1164 478144 1176
rect 478196 1164 478202 1216
rect 480898 1164 480904 1216
rect 480956 1204 480962 1216
rect 486418 1204 486424 1216
rect 480956 1176 486424 1204
rect 480956 1164 480962 1176
rect 486418 1164 486424 1176
rect 486476 1164 486482 1216
rect 486694 1164 486700 1216
rect 486752 1204 486758 1216
rect 492306 1204 492312 1216
rect 486752 1176 492312 1204
rect 486752 1164 486758 1176
rect 492306 1164 492312 1176
rect 492364 1164 492370 1216
rect 493594 1164 493600 1216
rect 493652 1204 493658 1216
rect 499390 1204 499396 1216
rect 493652 1176 499396 1204
rect 493652 1164 493658 1176
rect 499390 1164 499396 1176
rect 499448 1164 499454 1216
rect 500586 1164 500592 1216
rect 500644 1204 500650 1216
rect 506474 1204 506480 1216
rect 500644 1176 506480 1204
rect 500644 1164 500650 1176
rect 506474 1164 506480 1176
rect 506532 1164 506538 1216
rect 522666 1164 522672 1216
rect 522724 1204 522730 1216
rect 529014 1204 529020 1216
rect 522724 1176 529020 1204
rect 522724 1164 522730 1176
rect 529014 1164 529020 1176
rect 529072 1164 529078 1216
rect 530762 1164 530768 1216
rect 530820 1204 530826 1216
rect 537202 1204 537208 1216
rect 530820 1176 537208 1204
rect 530820 1164 530826 1176
rect 537202 1164 537208 1176
rect 537260 1164 537266 1216
rect 538858 1164 538864 1216
rect 538916 1204 538922 1216
rect 545482 1204 545488 1216
rect 538916 1176 545488 1204
rect 538916 1164 538922 1176
rect 545482 1164 545488 1176
rect 545540 1164 545546 1216
rect 550450 1164 550456 1216
rect 550508 1204 550514 1216
rect 557350 1204 557356 1216
rect 550508 1176 557356 1204
rect 550508 1164 550514 1176
rect 557350 1164 557356 1176
rect 557408 1164 557414 1216
rect 558454 1164 558460 1216
rect 558512 1204 558518 1216
rect 565630 1204 565636 1216
rect 558512 1176 565636 1204
rect 558512 1164 558518 1176
rect 565630 1164 565636 1176
rect 565688 1164 565694 1216
rect 569034 1164 569040 1216
rect 569092 1204 569098 1216
rect 576302 1204 576308 1216
rect 569092 1176 576308 1204
rect 569092 1164 569098 1176
rect 576302 1164 576308 1176
rect 576360 1164 576366 1216
rect 5626 1096 5632 1148
rect 5684 1136 5690 1148
rect 8662 1136 8668 1148
rect 5684 1108 8668 1136
rect 5684 1096 5690 1108
rect 8662 1096 8668 1108
rect 8720 1096 8726 1148
rect 111610 1096 111616 1148
rect 111668 1136 111674 1148
rect 113082 1136 113088 1148
rect 111668 1108 113088 1136
rect 111668 1096 111674 1108
rect 113082 1096 113088 1108
rect 113140 1096 113146 1148
rect 123478 1096 123484 1148
rect 123536 1136 123542 1148
rect 124766 1136 124772 1148
rect 123536 1108 124772 1136
rect 123536 1096 123542 1108
rect 124766 1096 124772 1108
rect 124824 1096 124830 1148
rect 320818 1096 320824 1148
rect 320876 1136 320882 1148
rect 323302 1136 323308 1148
rect 320876 1108 323308 1136
rect 320876 1096 320882 1108
rect 323302 1096 323308 1108
rect 323360 1096 323366 1148
rect 331122 1096 331128 1148
rect 331180 1136 331186 1148
rect 333882 1136 333888 1148
rect 331180 1108 333888 1136
rect 331180 1096 331186 1108
rect 333882 1096 333888 1108
rect 333940 1096 333946 1148
rect 360102 1096 360108 1148
rect 360160 1136 360166 1148
rect 363506 1136 363512 1148
rect 360160 1108 363512 1136
rect 360160 1096 360166 1108
rect 363506 1096 363512 1108
rect 363564 1096 363570 1148
rect 382182 1096 382188 1148
rect 382240 1136 382246 1148
rect 385954 1136 385960 1148
rect 382240 1108 385960 1136
rect 382240 1096 382246 1108
rect 385954 1096 385960 1108
rect 386012 1096 386018 1148
rect 389266 1096 389272 1148
rect 389324 1136 389330 1148
rect 393038 1136 393044 1148
rect 389324 1108 393044 1136
rect 389324 1096 389330 1108
rect 393038 1096 393044 1108
rect 393096 1096 393102 1148
rect 398466 1096 398472 1148
rect 398524 1136 398530 1148
rect 402514 1136 402520 1148
rect 398524 1108 402520 1136
rect 398524 1096 398530 1108
rect 402514 1096 402520 1108
rect 402572 1096 402578 1148
rect 404262 1096 404268 1148
rect 404320 1136 404326 1148
rect 408402 1136 408408 1148
rect 404320 1108 408408 1136
rect 404320 1096 404326 1108
rect 408402 1096 408408 1108
rect 408460 1096 408466 1148
rect 408954 1096 408960 1148
rect 409012 1136 409018 1148
rect 413094 1136 413100 1148
rect 409012 1108 413100 1136
rect 409012 1096 409018 1108
rect 413094 1096 413100 1108
rect 413152 1096 413158 1148
rect 415946 1096 415952 1148
rect 416004 1136 416010 1148
rect 420178 1136 420184 1148
rect 416004 1108 420184 1136
rect 416004 1096 416010 1108
rect 420178 1096 420184 1108
rect 420236 1096 420242 1148
rect 428642 1096 428648 1148
rect 428700 1136 428706 1148
rect 433242 1136 433248 1148
rect 428700 1108 433248 1136
rect 428700 1096 428706 1108
rect 433242 1096 433248 1108
rect 433300 1096 433306 1148
rect 439130 1096 439136 1148
rect 439188 1136 439194 1148
rect 443822 1136 443828 1148
rect 439188 1108 443828 1136
rect 439188 1096 439194 1108
rect 443822 1096 443828 1108
rect 443880 1096 443886 1148
rect 448422 1096 448428 1148
rect 448480 1136 448486 1148
rect 453298 1136 453304 1148
rect 448480 1108 453304 1136
rect 448480 1096 448486 1108
rect 453298 1096 453304 1108
rect 453356 1096 453362 1148
rect 454218 1096 454224 1148
rect 454276 1136 454282 1148
rect 459186 1136 459192 1148
rect 454276 1108 459192 1136
rect 454276 1096 454282 1108
rect 459186 1096 459192 1108
rect 459244 1096 459250 1148
rect 465810 1096 465816 1148
rect 465868 1136 465874 1148
rect 470686 1136 470692 1148
rect 465868 1108 470692 1136
rect 465868 1096 465874 1108
rect 470686 1096 470692 1108
rect 470744 1096 470750 1148
rect 482002 1096 482008 1148
rect 482060 1136 482066 1148
rect 487246 1136 487252 1148
rect 482060 1108 487252 1136
rect 482060 1096 482066 1108
rect 487246 1096 487252 1108
rect 487304 1096 487310 1148
rect 488994 1096 489000 1148
rect 489052 1136 489058 1148
rect 494698 1136 494704 1148
rect 489052 1108 494704 1136
rect 489052 1096 489058 1108
rect 494698 1096 494704 1108
rect 494756 1096 494762 1148
rect 501782 1096 501788 1148
rect 501840 1136 501846 1148
rect 507302 1136 507308 1148
rect 501840 1108 507308 1136
rect 501840 1096 501846 1108
rect 507302 1096 507308 1108
rect 507360 1096 507366 1148
rect 513282 1096 513288 1148
rect 513340 1136 513346 1148
rect 519538 1136 519544 1148
rect 513340 1108 519544 1136
rect 513340 1096 513346 1108
rect 519538 1096 519544 1108
rect 519596 1096 519602 1148
rect 523770 1096 523776 1148
rect 523828 1136 523834 1148
rect 530118 1136 530124 1148
rect 523828 1108 530124 1136
rect 523828 1096 523834 1108
rect 530118 1096 530124 1108
rect 530176 1096 530182 1148
rect 533062 1096 533068 1148
rect 533120 1136 533126 1148
rect 539594 1136 539600 1148
rect 533120 1108 539600 1136
rect 533120 1096 533126 1108
rect 539594 1096 539600 1108
rect 539652 1096 539658 1148
rect 543458 1096 543464 1148
rect 543516 1136 543522 1148
rect 550266 1136 550272 1148
rect 543516 1108 550272 1136
rect 543516 1096 543522 1108
rect 550266 1096 550272 1108
rect 550324 1096 550330 1148
rect 552750 1096 552756 1148
rect 552808 1136 552814 1148
rect 559742 1136 559748 1148
rect 552808 1108 559748 1136
rect 552808 1096 552814 1108
rect 559742 1096 559748 1108
rect 559800 1096 559806 1148
rect 567838 1096 567844 1148
rect 567896 1136 567902 1148
rect 575106 1136 575112 1148
rect 567896 1108 575112 1136
rect 567896 1096 567902 1108
rect 575106 1096 575112 1108
rect 575164 1096 575170 1148
rect 378778 1028 378784 1080
rect 378836 1068 378842 1080
rect 382366 1068 382372 1080
rect 378836 1040 382372 1068
rect 378836 1028 378842 1040
rect 382366 1028 382372 1040
rect 382424 1028 382430 1080
rect 386874 1028 386880 1080
rect 386932 1068 386938 1080
rect 390646 1068 390652 1080
rect 386932 1040 390652 1068
rect 386932 1028 386938 1040
rect 390646 1028 390652 1040
rect 390704 1028 390710 1080
rect 417050 1028 417056 1080
rect 417108 1068 417114 1080
rect 421374 1068 421380 1080
rect 417108 1040 421380 1068
rect 417108 1028 417114 1040
rect 421374 1028 421380 1040
rect 421432 1028 421438 1080
rect 437934 1028 437940 1080
rect 437992 1068 437998 1080
rect 442626 1068 442632 1080
rect 437992 1040 442632 1068
rect 437992 1028 437998 1040
rect 442626 1028 442632 1040
rect 442684 1028 442690 1080
rect 446030 1028 446036 1080
rect 446088 1068 446094 1080
rect 450906 1068 450912 1080
rect 446088 1040 450912 1068
rect 446088 1028 446094 1040
rect 450906 1028 450912 1040
rect 450964 1028 450970 1080
rect 455322 1028 455328 1080
rect 455380 1068 455386 1080
rect 460106 1068 460112 1080
rect 455380 1040 460112 1068
rect 455380 1028 455386 1040
rect 460106 1028 460112 1040
rect 460164 1028 460170 1080
rect 461118 1028 461124 1080
rect 461176 1068 461182 1080
rect 466270 1068 466276 1080
rect 461176 1040 466276 1068
rect 461176 1028 461182 1040
rect 466270 1028 466276 1040
rect 466328 1028 466334 1080
rect 466914 1028 466920 1080
rect 466972 1068 466978 1080
rect 472250 1068 472256 1080
rect 466972 1040 472256 1068
rect 466972 1028 466978 1040
rect 472250 1028 472256 1040
rect 472308 1028 472314 1080
rect 479702 1028 479708 1080
rect 479760 1068 479766 1080
rect 484854 1068 484860 1080
rect 479760 1040 484860 1068
rect 479760 1028 479766 1040
rect 484854 1028 484860 1040
rect 484912 1028 484918 1080
rect 491202 1028 491208 1080
rect 491260 1068 491266 1080
rect 497090 1068 497096 1080
rect 491260 1040 497096 1068
rect 491260 1028 491266 1040
rect 497090 1028 497096 1040
rect 497148 1028 497154 1080
rect 505186 1028 505192 1080
rect 505244 1068 505250 1080
rect 511258 1068 511264 1080
rect 505244 1040 511264 1068
rect 505244 1028 505250 1040
rect 511258 1028 511264 1040
rect 511316 1028 511322 1080
rect 512178 1028 512184 1080
rect 512236 1068 512242 1080
rect 517974 1068 517980 1080
rect 512236 1040 517980 1068
rect 512236 1028 512242 1040
rect 517974 1028 517980 1040
rect 518032 1028 518038 1080
rect 520182 1028 520188 1080
rect 520240 1068 520246 1080
rect 526622 1068 526628 1080
rect 520240 1040 526628 1068
rect 520240 1028 520246 1040
rect 526622 1028 526628 1040
rect 526680 1028 526686 1080
rect 529566 1028 529572 1080
rect 529624 1068 529630 1080
rect 536098 1068 536104 1080
rect 529624 1040 536104 1068
rect 529624 1028 529630 1040
rect 536098 1028 536104 1040
rect 536156 1028 536162 1080
rect 545850 1028 545856 1080
rect 545908 1068 545914 1080
rect 552658 1068 552664 1080
rect 545908 1040 552664 1068
rect 545908 1028 545914 1040
rect 552658 1028 552664 1040
rect 552716 1028 552722 1080
rect 559650 1028 559656 1080
rect 559708 1068 559714 1080
rect 566826 1068 566832 1080
rect 559708 1040 566832 1068
rect 559708 1028 559714 1040
rect 566826 1028 566832 1040
rect 566884 1028 566890 1080
rect 325418 960 325424 1012
rect 325476 1000 325482 1012
rect 327994 1000 328000 1012
rect 325476 972 328000 1000
rect 325476 960 325482 972
rect 327994 960 328000 972
rect 328052 960 328058 1012
rect 374178 960 374184 1012
rect 374236 1000 374242 1012
rect 377674 1000 377680 1012
rect 374236 972 377680 1000
rect 374236 960 374242 972
rect 377674 960 377680 972
rect 377732 960 377738 1012
rect 379882 960 379888 1012
rect 379940 1000 379946 1012
rect 383562 1000 383568 1012
rect 379940 972 383568 1000
rect 379940 960 379946 972
rect 383562 960 383568 972
rect 383620 960 383626 1012
rect 414750 960 414756 1012
rect 414808 1000 414814 1012
rect 418982 1000 418988 1012
rect 414808 972 418988 1000
rect 414808 960 414814 972
rect 418982 960 418988 972
rect 419040 960 419046 1012
rect 424042 960 424048 1012
rect 424100 1000 424106 1012
rect 428458 1000 428464 1012
rect 424100 972 428464 1000
rect 424100 960 424106 972
rect 428458 960 428464 972
rect 428516 960 428522 1012
rect 432138 960 432144 1012
rect 432196 1000 432202 1012
rect 436738 1000 436744 1012
rect 432196 972 436744 1000
rect 432196 960 432202 972
rect 436738 960 436744 972
rect 436796 960 436802 1012
rect 464614 960 464620 1012
rect 464672 1000 464678 1012
rect 469858 1000 469864 1012
rect 464672 972 469864 1000
rect 464672 960 464678 972
rect 469858 960 469864 972
rect 469916 960 469922 1012
rect 473906 960 473912 1012
rect 473964 1000 473970 1012
rect 479334 1000 479340 1012
rect 473964 972 479340 1000
rect 473964 960 473970 972
rect 479334 960 479340 972
rect 479392 960 479398 1012
rect 495986 960 495992 1012
rect 496044 1000 496050 1012
rect 501782 1000 501788 1012
rect 496044 972 501788 1000
rect 496044 960 496050 972
rect 501782 960 501788 972
rect 501840 960 501846 1012
rect 502886 960 502892 1012
rect 502944 1000 502950 1012
rect 508866 1000 508872 1012
rect 502944 972 508872 1000
rect 502944 960 502950 972
rect 508866 960 508872 972
rect 508924 960 508930 1012
rect 540054 960 540060 1012
rect 540112 1000 540118 1012
rect 546678 1000 546684 1012
rect 540112 972 546684 1000
rect 540112 960 540118 972
rect 546678 960 546684 972
rect 546736 960 546742 1012
rect 8754 892 8760 944
rect 8812 932 8818 944
rect 12158 932 12164 944
rect 8812 904 12164 932
rect 8812 892 8818 904
rect 12158 892 12164 904
rect 12216 892 12222 944
rect 121086 892 121092 944
rect 121144 932 121150 944
rect 122374 932 122380 944
rect 121144 904 122380 932
rect 121144 892 121150 904
rect 122374 892 122380 904
rect 122432 892 122438 944
rect 434346 892 434352 944
rect 434404 932 434410 944
rect 439130 932 439136 944
rect 434404 904 439136 932
rect 434404 892 434410 904
rect 439130 892 439136 904
rect 439188 892 439194 944
rect 463418 892 463424 944
rect 463476 932 463482 944
rect 468662 932 468668 944
rect 463476 904 468668 932
rect 463476 892 463482 904
rect 468662 892 468668 904
rect 468720 892 468726 944
rect 484302 892 484308 944
rect 484360 932 484366 944
rect 489914 932 489920 944
rect 484360 904 489920 932
rect 484360 892 484366 904
rect 489914 892 489920 904
rect 489972 892 489978 944
rect 347498 824 347504 876
rect 347556 864 347562 876
rect 350442 864 350448 876
rect 347556 836 350448 864
rect 347556 824 347562 836
rect 350442 824 350448 836
rect 350500 824 350506 876
rect 361390 824 361396 876
rect 361448 864 361454 876
rect 364610 864 364616 876
rect 361448 836 364616 864
rect 361448 824 361454 836
rect 364610 824 364616 836
rect 364668 824 364674 876
rect 368382 824 368388 876
rect 368440 864 368446 876
rect 371694 864 371700 876
rect 368440 836 371700 864
rect 368440 824 368446 836
rect 371694 824 371700 836
rect 371752 824 371758 876
rect 371786 824 371792 876
rect 371844 864 371850 876
rect 375282 864 375288 876
rect 371844 836 375288 864
rect 371844 824 371850 836
rect 375282 824 375288 836
rect 375340 824 375346 876
rect 384574 824 384580 876
rect 384632 864 384638 876
rect 388254 864 388260 876
rect 384632 836 388260 864
rect 384632 824 384638 836
rect 388254 824 388260 836
rect 388312 824 388318 876
rect 391566 824 391572 876
rect 391624 864 391630 876
rect 395338 864 395344 876
rect 391624 836 395344 864
rect 391624 824 391630 836
rect 395338 824 395344 836
rect 395396 824 395402 876
rect 397362 824 397368 876
rect 397420 864 397426 876
rect 401318 864 401324 876
rect 397420 836 401324 864
rect 397420 824 397426 836
rect 401318 824 401324 836
rect 401376 824 401382 876
rect 406654 824 406660 876
rect 406712 864 406718 876
rect 410794 864 410800 876
rect 406712 836 410800 864
rect 406712 824 406718 836
rect 410794 824 410800 836
rect 410852 824 410858 876
rect 419350 824 419356 876
rect 419408 864 419414 876
rect 423398 864 423404 876
rect 419408 836 423404 864
rect 419408 824 419414 836
rect 423398 824 423404 836
rect 423456 824 423462 876
rect 429838 824 429844 876
rect 429896 864 429902 876
rect 434438 864 434444 876
rect 429896 836 434444 864
rect 429896 824 429902 836
rect 434438 824 434444 836
rect 434496 824 434502 876
rect 443730 824 443736 876
rect 443788 864 443794 876
rect 448238 864 448244 876
rect 443788 836 448244 864
rect 443788 824 443794 836
rect 448238 824 448244 836
rect 448296 824 448302 876
rect 451826 824 451832 876
rect 451884 864 451890 876
rect 456518 864 456524 876
rect 451884 836 456524 864
rect 451884 824 451890 836
rect 456518 824 456524 836
rect 456576 824 456582 876
rect 476206 824 476212 876
rect 476264 864 476270 876
rect 481358 864 481364 876
rect 476264 836 481364 864
rect 476264 824 476270 836
rect 481358 824 481364 836
rect 481416 824 481422 876
rect 514478 824 514484 876
rect 514536 864 514542 876
rect 520734 864 520740 876
rect 514536 836 520740 864
rect 514536 824 514542 836
rect 520734 824 520740 836
rect 520792 824 520798 876
rect 521470 824 521476 876
rect 521528 864 521534 876
rect 527818 864 527824 876
rect 521528 836 527824 864
rect 521528 824 521534 836
rect 527818 824 527824 836
rect 527876 824 527882 876
rect 52546 688 52552 740
rect 52604 728 52610 740
rect 55030 728 55036 740
rect 52604 700 55036 728
rect 52604 688 52610 700
rect 55030 688 55036 700
rect 55088 688 55094 740
rect 59630 688 59636 740
rect 59688 728 59694 740
rect 61930 728 61936 740
rect 59688 700 61936 728
rect 59688 688 59694 700
rect 61930 688 61936 700
rect 61988 688 61994 740
rect 105722 688 105728 740
rect 105780 728 105786 740
rect 107286 728 107292 740
rect 105780 700 107292 728
rect 105780 688 105786 700
rect 107286 688 107292 700
rect 107344 688 107350 740
rect 274358 688 274364 740
rect 274416 728 274422 740
rect 276014 728 276020 740
rect 274416 700 276020 728
rect 274416 688 274422 700
rect 276014 688 276020 700
rect 276072 688 276078 740
rect 333514 688 333520 740
rect 333572 728 333578 740
rect 336274 728 336280 740
rect 333572 700 336280 728
rect 333572 688 333578 700
rect 336274 688 336280 700
rect 336332 688 336338 740
rect 338206 688 338212 740
rect 338264 728 338270 740
rect 340966 728 340972 740
rect 338264 700 340972 728
rect 338264 688 338270 700
rect 340966 688 340972 700
rect 341024 688 341030 740
rect 342806 688 342812 740
rect 342864 728 342870 740
rect 345750 728 345756 740
rect 342864 700 345756 728
rect 342864 688 342870 700
rect 345750 688 345756 700
rect 345808 688 345814 740
rect 346302 688 346308 740
rect 346360 728 346366 740
rect 349246 728 349252 740
rect 346360 700 349252 728
rect 346360 688 346366 700
rect 349246 688 349252 700
rect 349304 688 349310 740
rect 350902 688 350908 740
rect 350960 728 350966 740
rect 354030 728 354036 740
rect 350960 700 354036 728
rect 350960 688 350966 700
rect 354030 688 354036 700
rect 354088 688 354094 740
rect 365990 688 365996 740
rect 366048 728 366054 740
rect 369394 728 369400 740
rect 366048 700 369400 728
rect 366048 688 366054 700
rect 369394 688 369400 700
rect 369452 688 369458 740
rect 369486 688 369492 740
rect 369544 728 369550 740
rect 372890 728 372896 740
rect 369544 700 372896 728
rect 369544 688 369550 700
rect 372890 688 372896 700
rect 372948 688 372954 740
rect 544654 688 544660 740
rect 544712 728 544718 740
rect 551462 728 551468 740
rect 544712 700 551468 728
rect 544712 688 544718 700
rect 551462 688 551468 700
rect 551520 688 551526 740
rect 555142 688 555148 740
rect 555200 728 555206 740
rect 562042 728 562048 740
rect 555200 700 562048 728
rect 555200 688 555206 700
rect 562042 688 562048 700
rect 562100 688 562106 740
rect 494790 620 494796 672
rect 494848 660 494854 672
rect 500586 660 500592 672
rect 494848 632 500592 660
rect 494848 620 494854 632
rect 500586 620 500592 632
rect 500644 620 500650 672
rect 556246 620 556252 672
rect 556304 660 556310 672
rect 563146 660 563152 672
rect 556304 632 563152 660
rect 556304 620 556310 632
rect 563146 620 563152 632
rect 563204 620 563210 672
rect 69106 552 69112 604
rect 69164 592 69170 604
rect 71314 592 71320 604
rect 69164 564 71320 592
rect 69164 552 69170 564
rect 71314 552 71320 564
rect 71372 552 71378 604
rect 290642 552 290648 604
rect 290700 592 290706 604
rect 292574 592 292580 604
rect 290700 564 292580 592
rect 290700 552 290706 564
rect 292574 552 292580 564
rect 292632 552 292638 604
rect 304534 552 304540 604
rect 304592 592 304598 604
rect 306742 592 306748 604
rect 304592 564 306748 592
rect 304592 552 304598 564
rect 306742 552 306748 564
rect 306800 552 306806 604
rect 324222 552 324228 604
rect 324280 592 324286 604
rect 326798 592 326804 604
rect 324280 564 326804 592
rect 324280 552 324286 564
rect 326798 552 326804 564
rect 326856 552 326862 604
rect 327718 552 327724 604
rect 327776 592 327782 604
rect 330386 592 330392 604
rect 327776 564 330392 592
rect 327776 552 327782 564
rect 330386 552 330392 564
rect 330444 552 330450 604
rect 531866 552 531872 604
rect 531924 592 531930 604
rect 538398 592 538404 604
rect 531924 564 538404 592
rect 531924 552 531930 564
rect 538398 552 538404 564
rect 538456 552 538462 604
rect 544378 552 544384 604
rect 544436 552 544442 604
rect 549346 552 549352 604
rect 549404 592 549410 604
rect 556154 592 556160 604
rect 549404 564 556160 592
rect 549404 552 549410 564
rect 556154 552 556160 564
rect 556212 552 556218 604
rect 563330 552 563336 604
rect 563388 592 563394 604
rect 570322 592 570328 604
rect 563388 564 570328 592
rect 563388 552 563394 564
rect 570322 552 570328 564
rect 570380 552 570386 604
rect 537662 484 537668 536
rect 537720 524 537726 536
rect 544396 524 544424 552
rect 537720 496 544424 524
rect 537720 484 537726 496
rect 557534 484 557540 536
rect 557592 524 557598 536
rect 564618 524 564624 536
rect 557592 496 564624 524
rect 557592 484 557598 496
rect 564618 484 564624 496
rect 564676 484 564682 536
rect 535362 416 535368 468
rect 535420 456 535426 468
rect 542170 456 542176 468
rect 535420 428 542176 456
rect 535420 416 535426 428
rect 542170 416 542176 428
rect 542228 416 542234 468
rect 566642 416 566648 468
rect 566700 456 566706 468
rect 573726 456 573732 468
rect 566700 428 573732 456
rect 566700 416 566706 428
rect 573726 416 573732 428
rect 573784 416 573790 468
rect 383378 280 383384 332
rect 383436 320 383442 332
rect 386782 320 386788 332
rect 383436 292 386788 320
rect 383436 280 383442 292
rect 386782 280 386788 292
rect 386840 280 386846 332
rect 565446 280 565452 332
rect 565504 320 565510 332
rect 572898 320 572904 332
rect 565504 292 572904 320
rect 565504 280 565510 292
rect 572898 280 572904 292
rect 572956 280 572962 332
rect 576118 280 576124 332
rect 576176 320 576182 332
rect 583570 320 583576 332
rect 576176 292 583576 320
rect 576176 280 576182 292
rect 583570 280 583576 292
rect 583628 280 583634 332
rect 469306 212 469312 264
rect 469364 252 469370 264
rect 474182 252 474188 264
rect 469364 224 474188 252
rect 469364 212 469370 224
rect 474182 212 474188 224
rect 474240 212 474246 264
rect 508682 212 508688 264
rect 508740 252 508746 264
rect 514938 252 514944 264
rect 508740 224 514944 252
rect 508740 212 508746 224
rect 514938 212 514944 224
rect 514996 212 515002 264
rect 516778 212 516784 264
rect 516836 252 516842 264
rect 523218 252 523224 264
rect 516836 224 523224 252
rect 516836 212 516842 224
rect 523218 212 523224 224
rect 523276 212 523282 264
rect 553946 212 553952 264
rect 554004 252 554010 264
rect 560478 252 560484 264
rect 554004 224 560484 252
rect 554004 212 554010 224
rect 560478 212 560484 224
rect 560536 212 560542 264
rect 564250 212 564256 264
rect 564308 252 564314 264
rect 571334 252 571340 264
rect 564308 224 571340 252
rect 564308 212 564314 224
rect 571334 212 571340 224
rect 571392 212 571398 264
rect 574830 212 574836 264
rect 574888 252 574894 264
rect 581822 252 581828 264
rect 574888 224 581828 252
rect 574888 212 574894 224
rect 581822 212 581828 224
rect 581880 212 581886 264
rect 412450 144 412456 196
rect 412508 184 412514 196
rect 416866 184 416872 196
rect 412508 156 416872 184
rect 412508 144 412514 156
rect 416866 144 416872 156
rect 416924 144 416930 196
rect 470410 144 470416 196
rect 470468 184 470474 196
rect 475930 184 475936 196
rect 470468 156 475936 184
rect 470468 144 470474 156
rect 475930 144 475936 156
rect 475988 144 475994 196
rect 507486 144 507492 196
rect 507544 184 507550 196
rect 513374 184 513380 196
rect 507544 156 513380 184
rect 507544 144 507550 156
rect 513374 144 513380 156
rect 513432 144 513438 196
rect 392670 76 392676 128
rect 392728 116 392734 128
rect 396166 116 396172 128
rect 392728 88 396172 116
rect 392728 76 392734 88
rect 396166 76 396172 88
rect 396224 76 396230 128
rect 401962 76 401968 128
rect 402020 116 402026 128
rect 406194 116 406200 128
rect 402020 88 406200 116
rect 402020 76 402026 88
rect 406194 76 406200 88
rect 406252 76 406258 128
rect 421742 76 421748 128
rect 421800 116 421806 128
rect 425790 116 425796 128
rect 421800 88 425796 116
rect 421800 76 421806 88
rect 425790 76 425796 88
rect 425848 76 425854 128
rect 431034 76 431040 128
rect 431092 116 431098 128
rect 435174 116 435180 128
rect 431092 88 435180 116
rect 431092 76 431098 88
rect 435174 76 435180 88
rect 435232 76 435238 128
rect 460014 76 460020 128
rect 460072 116 460078 128
rect 464982 116 464988 128
rect 460072 88 464988 116
rect 460072 76 460078 88
rect 464982 76 464988 88
rect 465040 76 465046 128
rect 515674 76 515680 128
rect 515732 116 515738 128
rect 521654 116 521660 128
rect 515732 88 521660 116
rect 515732 76 515738 88
rect 521654 76 521660 88
rect 521712 76 521718 128
rect 524966 76 524972 128
rect 525024 116 525030 128
rect 531498 116 531504 128
rect 525024 88 531504 116
rect 525024 76 525030 88
rect 531498 76 531504 88
rect 531556 76 531562 128
rect 573634 76 573640 128
rect 573692 116 573698 128
rect 581178 116 581184 128
rect 573692 88 581184 116
rect 573692 76 573698 88
rect 581178 76 581184 88
rect 581236 76 581242 128
rect 354398 8 354404 60
rect 354456 48 354462 60
rect 357342 48 357348 60
rect 354456 20 357348 48
rect 354456 8 354462 20
rect 357342 8 357348 20
rect 357400 8 357406 60
rect 499206 8 499212 60
rect 499264 48 499270 60
rect 505554 48 505560 60
rect 499264 20 505560 48
rect 499264 8 499270 20
rect 505554 8 505560 20
rect 505612 8 505618 60
rect 506290 8 506296 60
rect 506348 48 506354 60
rect 512086 48 512092 60
rect 506348 20 512092 48
rect 506348 8 506354 20
rect 512086 8 512092 20
rect 512144 8 512150 60
rect 528462 8 528468 60
rect 528520 48 528526 60
rect 534534 48 534540 60
rect 528520 20 534540 48
rect 528520 8 528526 20
rect 534534 8 534540 20
rect 534592 8 534598 60
rect 536558 8 536564 60
rect 536616 48 536622 60
rect 542814 48 542820 60
rect 536616 20 542820 48
rect 536616 8 536622 20
rect 542814 8 542820 20
rect 542872 8 542878 60
rect 546954 8 546960 60
rect 547012 48 547018 60
rect 553946 48 553952 60
rect 547012 20 553952 48
rect 547012 8 547018 20
rect 553946 8 553952 20
rect 554004 8 554010 60
rect 572530 8 572536 60
rect 572588 48 572594 60
rect 579614 48 579620 60
rect 572588 20 579620 48
rect 572588 8 572594 20
rect 579614 8 579620 20
rect 579672 8 579678 60
<< via1 >>
rect 3884 700748 3936 700800
rect 8116 700748 8168 700800
rect 102048 700748 102100 700800
rect 105452 700748 105504 700800
rect 200028 700748 200080 700800
rect 202788 700748 202840 700800
rect 314476 700748 314528 700800
rect 316316 700748 316368 700800
rect 363512 700408 363564 700460
rect 364984 700408 365036 700460
rect 412456 700408 412508 700460
rect 413652 700408 413704 700460
rect 20352 700204 20404 700256
rect 24308 700204 24360 700256
rect 36728 700204 36780 700256
rect 40500 700204 40552 700256
rect 69388 700204 69440 700256
rect 72976 700204 73028 700256
rect 85764 700204 85816 700256
rect 89168 700204 89220 700256
rect 134708 700204 134760 700256
rect 137836 700204 137888 700256
rect 167368 700204 167420 700256
rect 170312 700204 170364 700256
rect 183744 700204 183796 700256
rect 186504 700204 186556 700256
rect 232780 700204 232832 700256
rect 235172 700204 235224 700256
rect 249064 700204 249116 700256
rect 251456 700204 251508 700256
rect 265440 700204 265492 700256
rect 267648 700204 267700 700256
rect 281816 700204 281868 700256
rect 283840 700204 283892 700256
rect 330760 700204 330812 700256
rect 332508 700204 332560 700256
rect 347136 700204 347188 700256
rect 348792 700204 348844 700256
rect 396172 700204 396224 700256
rect 397460 700204 397512 700256
rect 428832 700204 428884 700256
rect 429844 700204 429896 700256
rect 445208 700204 445260 700256
rect 446128 700204 446180 700256
rect 461492 700204 461544 700256
rect 462320 700204 462372 700256
rect 118424 700136 118476 700188
rect 121644 700136 121696 700188
rect 151084 700136 151136 700188
rect 154120 700136 154172 700188
rect 216404 700136 216456 700188
rect 218980 700136 219032 700188
rect 298008 700136 298060 700188
rect 300124 700136 300176 700188
rect 477868 700136 477920 700188
rect 478512 700136 478564 700188
rect 494244 700136 494296 700188
rect 494796 700136 494848 700188
rect 53012 700000 53064 700052
rect 56784 700000 56836 700052
rect 379796 699864 379848 699916
rect 381176 699864 381228 699916
rect 578332 644512 578384 644564
rect 580908 644512 580960 644564
rect 578884 257796 578936 257848
rect 580908 257796 580960 257848
rect 578516 151444 578568 151496
rect 580908 151444 580960 151496
rect 578332 44956 578384 45008
rect 579988 44956 580040 45008
rect 11152 3884 11204 3936
rect 14508 3884 14560 3936
rect 14740 3884 14792 3936
rect 18004 3884 18056 3936
rect 20628 3884 20680 3936
rect 23800 3884 23852 3936
rect 24216 3884 24268 3936
rect 27296 3884 27348 3936
rect 27712 3884 27764 3936
rect 30700 3884 30752 3936
rect 32404 3884 32456 3936
rect 35392 3884 35444 3936
rect 38384 3884 38436 3936
rect 41188 3884 41240 3936
rect 43076 3884 43128 3936
rect 45788 3884 45840 3936
rect 46664 3884 46716 3936
rect 49284 3884 49336 3936
rect 50160 3884 50212 3936
rect 52780 3884 52832 3936
rect 56048 3884 56100 3936
rect 58576 3884 58628 3936
rect 72608 3884 72660 3936
rect 74860 3884 74912 3936
rect 247636 3884 247688 3936
rect 248604 3884 248656 3936
rect 285908 3884 285960 3936
rect 287796 3884 287848 3936
rect 1676 3816 1728 3868
rect 5216 3816 5268 3868
rect 13544 3816 13596 3868
rect 16808 3816 16860 3868
rect 19432 3816 19484 3868
rect 22604 3816 22656 3868
rect 23020 3816 23072 3868
rect 26100 3816 26152 3868
rect 26516 3816 26568 3868
rect 29596 3816 29648 3868
rect 30104 3816 30156 3868
rect 33092 3816 33144 3868
rect 33600 3816 33652 3868
rect 36588 3816 36640 3868
rect 37188 3816 37240 3868
rect 39992 3816 40044 3868
rect 41880 3816 41932 3868
rect 44684 3816 44736 3868
rect 45468 3816 45520 3868
rect 48180 3816 48232 3868
rect 48964 3816 49016 3868
rect 51584 3816 51636 3868
rect 53748 3816 53800 3868
rect 56276 3816 56328 3868
rect 57244 3816 57296 3868
rect 59772 3816 59824 3868
rect 71504 3816 71556 3868
rect 73664 3816 73716 3868
rect 78588 3816 78640 3868
rect 80656 3816 80708 3868
rect 80888 3816 80940 3868
rect 82956 3816 83008 3868
rect 87972 3816 88024 3868
rect 89948 3816 90000 3868
rect 96252 3816 96304 3868
rect 98044 3816 98096 3868
rect 244140 3816 244192 3868
rect 245200 3816 245252 3868
rect 256928 3816 256980 3868
rect 258264 3816 258316 3868
rect 259228 3816 259280 3868
rect 260656 3816 260708 3868
rect 261620 3816 261672 3868
rect 262956 3816 263008 3868
rect 263920 3816 263972 3868
rect 265348 3816 265400 3868
rect 268520 3816 268572 3868
rect 270040 3816 270092 3868
rect 270820 3816 270872 3868
rect 272432 3816 272484 3868
rect 275512 3816 275564 3868
rect 277124 3816 277176 3868
rect 277812 3816 277864 3868
rect 279516 3816 279568 3868
rect 284804 3816 284856 3868
rect 286600 3816 286652 3868
rect 292900 3816 292952 3868
rect 294880 3816 294932 3868
rect 299892 3816 299944 3868
rect 301964 3816 302016 3868
rect 306792 3816 306844 3868
rect 309048 3816 309100 3868
rect 572 3748 624 3800
rect 4112 3748 4164 3800
rect 7656 3748 7708 3800
rect 11012 3748 11064 3800
rect 12348 3748 12400 3800
rect 15704 3748 15756 3800
rect 15936 3748 15988 3800
rect 19108 3748 19160 3800
rect 21824 3748 21876 3800
rect 24904 3748 24956 3800
rect 25320 3748 25372 3800
rect 28400 3748 28452 3800
rect 31300 3748 31352 3800
rect 34196 3748 34248 3800
rect 34796 3748 34848 3800
rect 37692 3748 37744 3800
rect 40684 3748 40736 3800
rect 43488 3748 43540 3800
rect 44272 3748 44324 3800
rect 46984 3748 47036 3800
rect 47860 3748 47912 3800
rect 50480 3748 50532 3800
rect 51356 3748 51408 3800
rect 53976 3748 54028 3800
rect 54944 3748 54996 3800
rect 57380 3748 57432 3800
rect 58440 3748 58492 3800
rect 60876 3748 60928 3800
rect 64328 3748 64380 3800
rect 66672 3748 66724 3800
rect 67088 3748 67140 3800
rect 69064 3748 69116 3800
rect 70308 3748 70360 3800
rect 72468 3748 72520 3800
rect 73804 3748 73856 3800
rect 75964 3748 76016 3800
rect 79692 3748 79744 3800
rect 81760 3748 81812 3800
rect 86868 3748 86920 3800
rect 88752 3748 88804 3800
rect 95148 3748 95200 3800
rect 96848 3748 96900 3800
rect 103336 3748 103388 3800
rect 104944 3748 104996 3800
rect 216356 3748 216408 3800
rect 216864 3748 216916 3800
rect 222152 3748 222204 3800
rect 222752 3748 222804 3800
rect 224452 3748 224504 3800
rect 225144 3748 225196 3800
rect 230248 3748 230300 3800
rect 231032 3748 231084 3800
rect 231444 3748 231496 3800
rect 232228 3748 232280 3800
rect 232548 3748 232600 3800
rect 233424 3748 233476 3800
rect 233744 3748 233796 3800
rect 234620 3748 234672 3800
rect 237240 3748 237292 3800
rect 238116 3748 238168 3800
rect 238344 3748 238396 3800
rect 239312 3748 239364 3800
rect 239540 3748 239592 3800
rect 240508 3748 240560 3800
rect 240736 3748 240788 3800
rect 241704 3748 241756 3800
rect 241840 3748 241892 3800
rect 242900 3748 242952 3800
rect 245336 3748 245388 3800
rect 246396 3748 246448 3800
rect 246532 3748 246584 3800
rect 247592 3748 247644 3800
rect 250028 3748 250080 3800
rect 251180 3748 251232 3800
rect 252328 3748 252380 3800
rect 253480 3748 253532 3800
rect 255824 3748 255876 3800
rect 257068 3748 257120 3800
rect 258124 3748 258176 3800
rect 259460 3748 259512 3800
rect 260424 3748 260476 3800
rect 261760 3748 261812 3800
rect 262724 3748 262776 3800
rect 264152 3748 264204 3800
rect 265024 3748 265076 3800
rect 266544 3748 266596 3800
rect 267416 3748 267468 3800
rect 268844 3748 268896 3800
rect 269716 3748 269768 3800
rect 271236 3748 271288 3800
rect 272016 3748 272068 3800
rect 273628 3748 273680 3800
rect 276708 3748 276760 3800
rect 278320 3748 278372 3800
rect 279008 3748 279060 3800
rect 280712 3748 280764 3800
rect 283608 3748 283660 3800
rect 285404 3748 285456 3800
rect 287104 3748 287156 3800
rect 288992 3748 289044 3800
rect 291704 3748 291756 3800
rect 293684 3748 293736 3800
rect 294096 3748 294148 3800
rect 296076 3748 296128 3800
rect 298696 3748 298748 3800
rect 300768 3748 300820 3800
rect 300996 3748 301048 3800
rect 303160 3748 303212 3800
rect 307988 3748 308040 3800
rect 310244 3748 310296 3800
rect 316084 3748 316136 3800
rect 318524 3748 318576 3800
rect 323076 3748 323128 3800
rect 325608 3748 325660 3800
rect 63224 3000 63276 3052
rect 65524 3000 65576 3052
rect 4068 2864 4120 2916
rect 7472 2864 7524 2916
rect 18236 2864 18288 2916
rect 21456 2864 21508 2916
rect 253388 2864 253440 2916
rect 254676 2864 254728 2916
rect 6460 2796 6512 2848
rect 9864 2796 9916 2848
rect 9956 2796 10008 2848
rect 13268 2796 13320 2848
rect 17040 2796 17092 2848
rect 20260 2796 20312 2848
rect 28908 2796 28960 2848
rect 31852 2796 31904 2848
rect 35992 2796 36044 2848
rect 38844 2796 38896 2848
rect 39580 2796 39632 2848
rect 42340 2796 42392 2848
rect 62028 2796 62080 2848
rect 64420 2796 64472 2848
rect 65524 2796 65576 2848
rect 67824 2796 67876 2848
rect 248880 2796 248932 2848
rect 249984 2796 250036 2848
rect 251088 2796 251140 2848
rect 252376 2796 252428 2848
rect 254584 2796 254636 2848
rect 255872 2796 255924 2848
rect 309232 2796 309284 2848
rect 311440 2796 311492 2848
rect 315028 2796 315080 2848
rect 317328 2796 317380 2848
rect 411168 2796 411220 2848
rect 415492 2796 415544 2848
rect 440148 2796 440200 2848
rect 445024 2796 445076 2848
rect 449532 2796 449584 2848
rect 454500 2796 454552 2848
rect 478512 2796 478564 2848
rect 484032 2796 484084 2848
rect 487804 2796 487856 2848
rect 493508 2796 493560 2848
rect 3240 1300 3292 1352
rect 6368 1300 6420 1352
rect 60832 1300 60884 1352
rect 63316 1300 63368 1352
rect 67916 1300 67968 1352
rect 70124 1300 70176 1352
rect 76196 1300 76248 1352
rect 78220 1300 78272 1352
rect 83280 1300 83332 1352
rect 85212 1300 85264 1352
rect 85672 1300 85724 1352
rect 87512 1300 87564 1352
rect 89168 1300 89220 1352
rect 91008 1300 91060 1352
rect 91560 1300 91612 1352
rect 93308 1300 93360 1352
rect 93952 1300 94004 1352
rect 95700 1300 95752 1352
rect 97448 1300 97500 1352
rect 99104 1300 99156 1352
rect 101036 1300 101088 1352
rect 102600 1300 102652 1352
rect 104532 1300 104584 1352
rect 106096 1300 106148 1352
rect 106924 1300 106976 1352
rect 108396 1300 108448 1352
rect 109316 1300 109368 1352
rect 110696 1300 110748 1352
rect 112812 1300 112864 1352
rect 114192 1300 114244 1352
rect 116400 1300 116452 1352
rect 117688 1300 117740 1352
rect 119896 1300 119948 1352
rect 121184 1300 121236 1352
rect 125876 1300 125928 1352
rect 126980 1300 127032 1352
rect 129372 1300 129424 1352
rect 130476 1300 130528 1352
rect 130568 1300 130620 1352
rect 131580 1300 131632 1352
rect 131764 1300 131816 1352
rect 132776 1300 132828 1352
rect 132960 1300 133012 1352
rect 133972 1300 134024 1352
rect 137652 1300 137704 1352
rect 138572 1300 138624 1352
rect 144736 1300 144788 1352
rect 145564 1300 145616 1352
rect 145932 1300 145984 1352
rect 146668 1300 146720 1352
rect 148324 1300 148376 1352
rect 149060 1300 149112 1352
rect 154212 1300 154264 1352
rect 154856 1300 154908 1352
rect 162492 1300 162544 1352
rect 162952 1300 163004 1352
rect 266268 1300 266320 1352
rect 267740 1300 267792 1352
rect 273168 1300 273220 1352
rect 274824 1300 274876 1352
rect 280068 1300 280120 1352
rect 281908 1300 281960 1352
rect 282552 1300 282604 1352
rect 284300 1300 284352 1352
rect 288348 1300 288400 1352
rect 290188 1300 290240 1352
rect 295248 1300 295300 1352
rect 297272 1300 297324 1352
rect 297548 1300 297600 1352
rect 299664 1300 299716 1352
rect 302148 1300 302200 1352
rect 304356 1300 304408 1352
rect 305736 1300 305788 1352
rect 307944 1300 307996 1352
rect 310336 1300 310388 1352
rect 312636 1300 312688 1352
rect 313832 1300 313884 1352
rect 316224 1300 316276 1352
rect 317236 1300 317288 1352
rect 319720 1300 319772 1352
rect 321928 1300 321980 1352
rect 324412 1300 324464 1352
rect 326620 1300 326672 1352
rect 329196 1300 329248 1352
rect 332416 1300 332468 1352
rect 335084 1300 335136 1352
rect 335912 1300 335964 1352
rect 338672 1300 338724 1352
rect 339316 1300 339368 1352
rect 342168 1300 342220 1352
rect 345112 1300 345164 1352
rect 348056 1300 348108 1352
rect 349804 1300 349856 1352
rect 352840 1300 352892 1352
rect 353208 1300 353260 1352
rect 356336 1300 356388 1352
rect 356704 1300 356756 1352
rect 359924 1300 359976 1352
rect 362592 1300 362644 1352
rect 365812 1300 365864 1352
rect 367192 1300 367244 1352
rect 370596 1300 370648 1352
rect 370688 1300 370740 1352
rect 374092 1300 374144 1352
rect 376392 1300 376444 1352
rect 379980 1300 380032 1352
rect 385776 1300 385828 1352
rect 389456 1300 389508 1352
rect 395068 1300 395120 1352
rect 398932 1300 398984 1352
rect 399668 1300 399720 1352
rect 403624 1300 403676 1352
rect 405464 1300 405516 1352
rect 409604 1300 409656 1352
rect 413560 1300 413612 1352
rect 417884 1300 417936 1352
rect 422852 1300 422904 1352
rect 427268 1300 427320 1352
rect 427544 1300 427596 1352
rect 431868 1300 431920 1352
rect 433248 1300 433300 1352
rect 437848 1300 437900 1352
rect 441436 1300 441488 1352
rect 445852 1300 445904 1352
rect 447232 1300 447284 1352
rect 452108 1300 452160 1352
rect 453028 1300 453080 1352
rect 458088 1300 458140 1352
rect 458824 1300 458876 1352
rect 463976 1300 464028 1352
rect 471612 1300 471664 1352
rect 476580 1300 476632 1352
rect 477408 1300 477460 1352
rect 482468 1300 482520 1352
rect 483204 1300 483256 1352
rect 488816 1300 488868 1352
rect 490104 1300 490156 1352
rect 495532 1300 495584 1352
rect 497096 1300 497148 1352
rect 502984 1300 503036 1352
rect 504088 1300 504140 1352
rect 509700 1300 509752 1352
rect 509884 1300 509936 1352
rect 515772 1300 515824 1352
rect 519176 1300 519228 1352
rect 525432 1300 525484 1352
rect 526076 1300 526128 1352
rect 532148 1300 532200 1352
rect 534264 1300 534316 1352
rect 540428 1300 540480 1352
rect 542268 1300 542320 1352
rect 549076 1300 549128 1352
rect 551652 1300 551704 1352
rect 558552 1300 558604 1352
rect 560944 1300 560996 1352
rect 568028 1300 568080 1352
rect 571248 1300 571300 1352
rect 578608 1300 578660 1352
rect 75000 1232 75052 1284
rect 77116 1232 77168 1284
rect 77392 1232 77444 1284
rect 79416 1232 79468 1284
rect 82084 1232 82136 1284
rect 84016 1232 84068 1284
rect 84476 1232 84528 1284
rect 86408 1232 86460 1284
rect 90364 1232 90416 1284
rect 92204 1232 92256 1284
rect 92756 1232 92808 1284
rect 94504 1232 94556 1284
rect 98644 1232 98696 1284
rect 100300 1232 100352 1284
rect 102232 1232 102284 1284
rect 103796 1232 103848 1284
rect 108120 1232 108172 1284
rect 109592 1232 109644 1284
rect 110512 1232 110564 1284
rect 111892 1232 111944 1284
rect 115204 1232 115256 1284
rect 116584 1232 116636 1284
rect 117596 1232 117648 1284
rect 118884 1232 118936 1284
rect 122288 1232 122340 1284
rect 123484 1232 123536 1284
rect 124680 1232 124732 1284
rect 125784 1232 125836 1284
rect 128176 1232 128228 1284
rect 129280 1232 129332 1284
rect 136456 1232 136508 1284
rect 137376 1232 137428 1284
rect 138848 1232 138900 1284
rect 139768 1232 139820 1284
rect 140044 1232 140096 1284
rect 140872 1232 140924 1284
rect 281356 1232 281408 1284
rect 283104 1232 283156 1284
rect 289452 1232 289504 1284
rect 291384 1232 291436 1284
rect 296444 1232 296496 1284
rect 298468 1232 298520 1284
rect 303344 1232 303396 1284
rect 305552 1232 305604 1284
rect 312544 1232 312596 1284
rect 315028 1232 315080 1284
rect 318432 1232 318484 1284
rect 320916 1232 320968 1284
rect 328920 1232 328972 1284
rect 331588 1232 331640 1284
rect 334716 1232 334768 1284
rect 337476 1232 337528 1284
rect 340512 1232 340564 1284
rect 343364 1232 343416 1284
rect 344008 1232 344060 1284
rect 346952 1232 347004 1284
rect 348608 1232 348660 1284
rect 351644 1232 351696 1284
rect 352104 1232 352156 1284
rect 355232 1232 355284 1284
rect 355600 1232 355652 1284
rect 358728 1232 358780 1284
rect 359096 1232 359148 1284
rect 362316 1232 362368 1284
rect 363696 1232 363748 1284
rect 367008 1232 367060 1284
rect 372988 1232 373040 1284
rect 376484 1232 376536 1284
rect 377588 1232 377640 1284
rect 381176 1232 381228 1284
rect 388076 1232 388128 1284
rect 391848 1232 391900 1284
rect 393872 1232 393924 1284
rect 397736 1232 397788 1284
rect 403164 1232 403216 1284
rect 407212 1232 407264 1284
rect 410064 1232 410116 1284
rect 414296 1232 414348 1284
rect 418252 1232 418304 1284
rect 422576 1232 422628 1284
rect 426348 1232 426400 1284
rect 430856 1232 430908 1284
rect 435640 1232 435692 1284
rect 439964 1232 440016 1284
rect 442632 1232 442684 1284
rect 447416 1232 447468 1284
rect 457628 1232 457680 1284
rect 462412 1232 462464 1284
rect 468116 1232 468168 1284
rect 473084 1232 473136 1284
rect 475108 1232 475160 1284
rect 480536 1232 480588 1284
rect 485504 1232 485556 1284
rect 490748 1232 490800 1284
rect 492496 1232 492548 1284
rect 498200 1232 498252 1284
rect 498292 1232 498344 1284
rect 503812 1232 503864 1284
rect 510988 1232 511040 1284
rect 517152 1232 517204 1284
rect 517980 1232 518032 1284
rect 523868 1232 523920 1284
rect 527272 1232 527324 1284
rect 533712 1232 533764 1284
rect 541164 1232 541216 1284
rect 547880 1232 547932 1284
rect 548156 1232 548208 1284
rect 554964 1232 555016 1284
rect 562048 1232 562100 1284
rect 569132 1232 569184 1284
rect 570144 1232 570196 1284
rect 577412 1232 577464 1284
rect 99840 1164 99892 1216
rect 101496 1164 101548 1216
rect 114008 1164 114060 1216
rect 115388 1164 115440 1216
rect 311532 1164 311584 1216
rect 313832 1164 313884 1216
rect 319628 1164 319680 1216
rect 322112 1164 322164 1216
rect 330024 1164 330076 1216
rect 332692 1164 332744 1216
rect 337016 1164 337068 1216
rect 339868 1164 339920 1216
rect 341708 1164 341760 1216
rect 344560 1164 344612 1216
rect 357900 1164 357952 1216
rect 361120 1164 361172 1216
rect 364892 1164 364944 1216
rect 368204 1164 368256 1216
rect 375288 1164 375340 1216
rect 378876 1164 378928 1216
rect 381084 1164 381136 1216
rect 384764 1164 384816 1216
rect 390376 1164 390428 1216
rect 394240 1164 394292 1216
rect 396172 1164 396224 1216
rect 400128 1164 400180 1216
rect 400864 1164 400916 1216
rect 404820 1164 404872 1216
rect 407764 1164 407816 1216
rect 411904 1164 411956 1216
rect 420552 1164 420604 1216
rect 424968 1164 425020 1216
rect 425152 1164 425204 1216
rect 429660 1164 429712 1216
rect 436744 1164 436796 1216
rect 441528 1164 441580 1216
rect 444932 1164 444984 1216
rect 449808 1164 449860 1216
rect 450728 1164 450780 1216
rect 455696 1164 455748 1216
rect 456524 1164 456576 1216
rect 461584 1164 461636 1216
rect 462228 1164 462280 1216
rect 467472 1164 467524 1216
rect 472716 1164 472768 1216
rect 478144 1164 478196 1216
rect 480904 1164 480956 1216
rect 486424 1164 486476 1216
rect 486700 1164 486752 1216
rect 492312 1164 492364 1216
rect 493600 1164 493652 1216
rect 499396 1164 499448 1216
rect 500592 1164 500644 1216
rect 506480 1164 506532 1216
rect 522672 1164 522724 1216
rect 529020 1164 529072 1216
rect 530768 1164 530820 1216
rect 537208 1164 537260 1216
rect 538864 1164 538916 1216
rect 545488 1164 545540 1216
rect 550456 1164 550508 1216
rect 557356 1164 557408 1216
rect 558460 1164 558512 1216
rect 565636 1164 565688 1216
rect 569040 1164 569092 1216
rect 576308 1164 576360 1216
rect 5632 1096 5684 1148
rect 8668 1096 8720 1148
rect 111616 1096 111668 1148
rect 113088 1096 113140 1148
rect 123484 1096 123536 1148
rect 124772 1096 124824 1148
rect 320824 1096 320876 1148
rect 323308 1096 323360 1148
rect 331128 1096 331180 1148
rect 333888 1096 333940 1148
rect 360108 1096 360160 1148
rect 363512 1096 363564 1148
rect 382188 1096 382240 1148
rect 385960 1096 386012 1148
rect 389272 1096 389324 1148
rect 393044 1096 393096 1148
rect 398472 1096 398524 1148
rect 402520 1096 402572 1148
rect 404268 1096 404320 1148
rect 408408 1096 408460 1148
rect 408960 1096 409012 1148
rect 413100 1096 413152 1148
rect 415952 1096 416004 1148
rect 420184 1096 420236 1148
rect 428648 1096 428700 1148
rect 433248 1096 433300 1148
rect 439136 1096 439188 1148
rect 443828 1096 443880 1148
rect 448428 1096 448480 1148
rect 453304 1096 453356 1148
rect 454224 1096 454276 1148
rect 459192 1096 459244 1148
rect 465816 1096 465868 1148
rect 470692 1096 470744 1148
rect 482008 1096 482060 1148
rect 487252 1096 487304 1148
rect 489000 1096 489052 1148
rect 494704 1096 494756 1148
rect 501788 1096 501840 1148
rect 507308 1096 507360 1148
rect 513288 1096 513340 1148
rect 519544 1096 519596 1148
rect 523776 1096 523828 1148
rect 530124 1096 530176 1148
rect 533068 1096 533120 1148
rect 539600 1096 539652 1148
rect 543464 1096 543516 1148
rect 550272 1096 550324 1148
rect 552756 1096 552808 1148
rect 559748 1096 559800 1148
rect 567844 1096 567896 1148
rect 575112 1096 575164 1148
rect 378784 1028 378836 1080
rect 382372 1028 382424 1080
rect 386880 1028 386932 1080
rect 390652 1028 390704 1080
rect 417056 1028 417108 1080
rect 421380 1028 421432 1080
rect 437940 1028 437992 1080
rect 442632 1028 442684 1080
rect 446036 1028 446088 1080
rect 450912 1028 450964 1080
rect 455328 1028 455380 1080
rect 460112 1028 460164 1080
rect 461124 1028 461176 1080
rect 466276 1028 466328 1080
rect 466920 1028 466972 1080
rect 472256 1028 472308 1080
rect 479708 1028 479760 1080
rect 484860 1028 484912 1080
rect 491208 1028 491260 1080
rect 497096 1028 497148 1080
rect 505192 1028 505244 1080
rect 511264 1028 511316 1080
rect 512184 1028 512236 1080
rect 517980 1028 518032 1080
rect 520188 1028 520240 1080
rect 526628 1028 526680 1080
rect 529572 1028 529624 1080
rect 536104 1028 536156 1080
rect 545856 1028 545908 1080
rect 552664 1028 552716 1080
rect 559656 1028 559708 1080
rect 566832 1028 566884 1080
rect 325424 960 325476 1012
rect 328000 960 328052 1012
rect 374184 960 374236 1012
rect 377680 960 377732 1012
rect 379888 960 379940 1012
rect 383568 960 383620 1012
rect 414756 960 414808 1012
rect 418988 960 419040 1012
rect 424048 960 424100 1012
rect 428464 960 428516 1012
rect 432144 960 432196 1012
rect 436744 960 436796 1012
rect 464620 960 464672 1012
rect 469864 960 469916 1012
rect 473912 960 473964 1012
rect 479340 960 479392 1012
rect 495992 960 496044 1012
rect 501788 960 501840 1012
rect 502892 960 502944 1012
rect 508872 960 508924 1012
rect 540060 960 540112 1012
rect 546684 960 546736 1012
rect 8760 892 8812 944
rect 12164 892 12216 944
rect 121092 892 121144 944
rect 122380 892 122432 944
rect 434352 892 434404 944
rect 439136 892 439188 944
rect 463424 892 463476 944
rect 468668 892 468720 944
rect 484308 892 484360 944
rect 489920 892 489972 944
rect 347504 824 347556 876
rect 350448 824 350500 876
rect 361396 824 361448 876
rect 364616 824 364668 876
rect 368388 824 368440 876
rect 371700 824 371752 876
rect 371792 824 371844 876
rect 375288 824 375340 876
rect 384580 824 384632 876
rect 388260 824 388312 876
rect 391572 824 391624 876
rect 395344 824 395396 876
rect 397368 824 397420 876
rect 401324 824 401376 876
rect 406660 824 406712 876
rect 410800 824 410852 876
rect 419356 824 419408 876
rect 423404 824 423456 876
rect 429844 824 429896 876
rect 434444 824 434496 876
rect 443736 824 443788 876
rect 448244 824 448296 876
rect 451832 824 451884 876
rect 456524 824 456576 876
rect 476212 824 476264 876
rect 481364 824 481416 876
rect 514484 824 514536 876
rect 520740 824 520792 876
rect 521476 824 521528 876
rect 527824 824 527876 876
rect 52552 688 52604 740
rect 55036 688 55088 740
rect 59636 688 59688 740
rect 61936 688 61988 740
rect 105728 688 105780 740
rect 107292 688 107344 740
rect 274364 688 274416 740
rect 276020 688 276072 740
rect 333520 688 333572 740
rect 336280 688 336332 740
rect 338212 688 338264 740
rect 340972 688 341024 740
rect 342812 688 342864 740
rect 345756 688 345808 740
rect 346308 688 346360 740
rect 349252 688 349304 740
rect 350908 688 350960 740
rect 354036 688 354088 740
rect 365996 688 366048 740
rect 369400 688 369452 740
rect 369492 688 369544 740
rect 372896 688 372948 740
rect 544660 688 544712 740
rect 551468 688 551520 740
rect 555148 688 555200 740
rect 562048 688 562100 740
rect 494796 620 494848 672
rect 500592 620 500644 672
rect 556252 620 556304 672
rect 563152 620 563204 672
rect 69112 552 69164 604
rect 71320 552 71372 604
rect 290648 552 290700 604
rect 292580 552 292632 604
rect 304540 552 304592 604
rect 306748 552 306800 604
rect 324228 552 324280 604
rect 326804 552 326856 604
rect 327724 552 327776 604
rect 330392 552 330444 604
rect 531872 552 531924 604
rect 538404 552 538456 604
rect 544384 552 544436 604
rect 549352 552 549404 604
rect 556160 552 556212 604
rect 563336 552 563388 604
rect 570328 552 570380 604
rect 537668 484 537720 536
rect 557540 484 557592 536
rect 564624 484 564676 536
rect 535368 416 535420 468
rect 542176 416 542228 468
rect 566648 416 566700 468
rect 573732 416 573784 468
rect 383384 280 383436 332
rect 386788 280 386840 332
rect 565452 280 565504 332
rect 572904 280 572956 332
rect 576124 280 576176 332
rect 583576 280 583628 332
rect 469312 212 469364 264
rect 474188 212 474240 264
rect 508688 212 508740 264
rect 514944 212 514996 264
rect 516784 212 516836 264
rect 523224 212 523276 264
rect 553952 212 554004 264
rect 560484 212 560536 264
rect 564256 212 564308 264
rect 571340 212 571392 264
rect 574836 212 574888 264
rect 581828 212 581880 264
rect 412456 144 412508 196
rect 416872 144 416924 196
rect 470416 144 470468 196
rect 475936 144 475988 196
rect 507492 144 507544 196
rect 513380 144 513432 196
rect 392676 76 392728 128
rect 396172 76 396224 128
rect 401968 76 402020 128
rect 406200 76 406252 128
rect 421748 76 421800 128
rect 425796 76 425848 128
rect 431040 76 431092 128
rect 435180 76 435232 128
rect 460020 76 460072 128
rect 464988 76 465040 128
rect 515680 76 515732 128
rect 521660 76 521712 128
rect 524972 76 525024 128
rect 531504 76 531556 128
rect 573640 76 573692 128
rect 581184 76 581236 128
rect 354404 8 354456 60
rect 357348 8 357400 60
rect 499212 8 499264 60
rect 505560 8 505612 60
rect 506296 8 506348 60
rect 512092 8 512144 60
rect 528468 8 528520 60
rect 534540 8 534592 60
rect 536564 8 536616 60
rect 542820 8 542872 60
rect 546960 8 547012 60
rect 553952 8 554004 60
rect 572536 8 572588 60
rect 579620 8 579672 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510632 703582 510844 703610
rect 8128 700806 8156 703520
rect 3884 700800 3936 700806
rect 3884 700742 3936 700748
rect 8116 700800 8168 700806
rect 8116 700742 8168 700748
rect 3514 697976 3570 697985
rect 3896 697966 3924 700742
rect 24320 700262 24348 703520
rect 40512 700262 40540 703520
rect 20352 700256 20404 700262
rect 20352 700198 20404 700204
rect 24308 700256 24360 700262
rect 24308 700198 24360 700204
rect 36728 700256 36780 700262
rect 36728 700198 36780 700204
rect 40500 700256 40552 700262
rect 40500 700198 40552 700204
rect 20364 698170 20392 700198
rect 36740 698170 36768 700198
rect 56796 700058 56824 703520
rect 72988 700262 73016 703520
rect 89180 700262 89208 703520
rect 105464 700806 105492 703520
rect 102048 700800 102100 700806
rect 102048 700742 102100 700748
rect 105452 700800 105504 700806
rect 105452 700742 105504 700748
rect 69388 700256 69440 700262
rect 69388 700198 69440 700204
rect 72976 700256 73028 700262
rect 72976 700198 73028 700204
rect 85764 700256 85816 700262
rect 85764 700198 85816 700204
rect 89168 700256 89220 700262
rect 89168 700198 89220 700204
rect 53012 700052 53064 700058
rect 53012 699994 53064 700000
rect 56784 700052 56836 700058
rect 56784 699994 56836 700000
rect 53024 698170 53052 699994
rect 69400 698170 69428 700198
rect 85776 698170 85804 700198
rect 102060 698170 102088 700742
rect 121656 700194 121684 703520
rect 137848 700262 137876 703520
rect 134708 700256 134760 700262
rect 134708 700198 134760 700204
rect 137836 700256 137888 700262
rect 137836 700198 137888 700204
rect 118424 700188 118476 700194
rect 118424 700130 118476 700136
rect 121644 700188 121696 700194
rect 121644 700130 121696 700136
rect 118436 698170 118464 700130
rect 134720 698170 134748 700198
rect 154132 700194 154160 703520
rect 170324 700262 170352 703520
rect 186516 700262 186544 703520
rect 202800 700806 202828 703520
rect 200028 700800 200080 700806
rect 200028 700742 200080 700748
rect 202788 700800 202840 700806
rect 202788 700742 202840 700748
rect 167368 700256 167420 700262
rect 167368 700198 167420 700204
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 183744 700256 183796 700262
rect 183744 700198 183796 700204
rect 186504 700256 186556 700262
rect 186504 700198 186556 700204
rect 151084 700188 151136 700194
rect 151084 700130 151136 700136
rect 154120 700188 154172 700194
rect 154120 700130 154172 700136
rect 151096 698170 151124 700130
rect 167380 698170 167408 700198
rect 183756 698170 183784 700198
rect 20316 698142 20392 698170
rect 36692 698142 36768 698170
rect 52976 698142 53052 698170
rect 69352 698142 69428 698170
rect 85728 698142 85804 698170
rect 102012 698142 102088 698170
rect 118388 698142 118464 698170
rect 134672 698142 134748 698170
rect 151048 698142 151124 698170
rect 167332 698142 167408 698170
rect 183708 698142 183784 698170
rect 200040 698170 200068 700742
rect 218992 700194 219020 703520
rect 235184 700262 235212 703520
rect 251468 700262 251496 703520
rect 267660 700262 267688 703520
rect 283852 700262 283880 703520
rect 232780 700256 232832 700262
rect 232780 700198 232832 700204
rect 235172 700256 235224 700262
rect 235172 700198 235224 700204
rect 249064 700256 249116 700262
rect 249064 700198 249116 700204
rect 251456 700256 251508 700262
rect 251456 700198 251508 700204
rect 265440 700256 265492 700262
rect 265440 700198 265492 700204
rect 267648 700256 267700 700262
rect 267648 700198 267700 700204
rect 281816 700256 281868 700262
rect 281816 700198 281868 700204
rect 283840 700256 283892 700262
rect 283840 700198 283892 700204
rect 216404 700188 216456 700194
rect 216404 700130 216456 700136
rect 218980 700188 219032 700194
rect 218980 700130 219032 700136
rect 216416 698170 216444 700130
rect 232792 698170 232820 700198
rect 249076 698170 249104 700198
rect 265452 698170 265480 700198
rect 281828 698170 281856 700198
rect 300136 700194 300164 703520
rect 316328 700806 316356 703520
rect 314476 700800 314528 700806
rect 314476 700742 314528 700748
rect 316316 700800 316368 700806
rect 316316 700742 316368 700748
rect 298008 700188 298060 700194
rect 298008 700130 298060 700136
rect 300124 700188 300176 700194
rect 300124 700130 300176 700136
rect 200040 698142 200112 698170
rect 3896 697938 4046 697966
rect 20316 697959 20344 698142
rect 36692 697959 36720 698142
rect 52976 697959 53004 698142
rect 69352 697959 69380 698142
rect 85728 697959 85756 698142
rect 102012 697959 102040 698142
rect 118388 697959 118416 698142
rect 134672 697959 134700 698142
rect 151048 697959 151076 698142
rect 167332 697959 167360 698142
rect 183708 697959 183736 698142
rect 200084 697959 200112 698142
rect 216368 698142 216444 698170
rect 232744 698142 232820 698170
rect 249028 698142 249104 698170
rect 265404 698142 265480 698170
rect 281780 698142 281856 698170
rect 298020 698170 298048 700130
rect 314488 698170 314516 700742
rect 332520 700262 332548 703520
rect 348804 700262 348832 703520
rect 364996 700466 365024 703520
rect 363512 700460 363564 700466
rect 363512 700402 363564 700408
rect 364984 700460 365036 700466
rect 364984 700402 365036 700408
rect 330760 700256 330812 700262
rect 330760 700198 330812 700204
rect 332508 700256 332560 700262
rect 332508 700198 332560 700204
rect 347136 700256 347188 700262
rect 347136 700198 347188 700204
rect 348792 700256 348844 700262
rect 348792 700198 348844 700204
rect 330772 698170 330800 700198
rect 347148 698170 347176 700198
rect 363524 698170 363552 700402
rect 381188 699922 381216 703520
rect 397472 700262 397500 703520
rect 413664 700466 413692 703520
rect 412456 700460 412508 700466
rect 412456 700402 412508 700408
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 396172 700256 396224 700262
rect 396172 700198 396224 700204
rect 397460 700256 397512 700262
rect 397460 700198 397512 700204
rect 379796 699916 379848 699922
rect 379796 699858 379848 699864
rect 381176 699916 381228 699922
rect 381176 699858 381228 699864
rect 379808 698170 379836 699858
rect 396184 698170 396212 700198
rect 412468 698170 412496 700402
rect 429856 700262 429884 703520
rect 446140 700262 446168 703520
rect 462332 700262 462360 703520
rect 428832 700256 428884 700262
rect 428832 700198 428884 700204
rect 429844 700256 429896 700262
rect 429844 700198 429896 700204
rect 445208 700256 445260 700262
rect 445208 700198 445260 700204
rect 446128 700256 446180 700262
rect 446128 700198 446180 700204
rect 461492 700256 461544 700262
rect 461492 700198 461544 700204
rect 462320 700256 462372 700262
rect 462320 700198 462372 700204
rect 428844 698170 428872 700198
rect 445220 698170 445248 700198
rect 461504 698170 461532 700198
rect 478524 700194 478552 703520
rect 494808 700194 494836 703520
rect 477868 700188 477920 700194
rect 477868 700130 477920 700136
rect 478512 700188 478564 700194
rect 478512 700130 478564 700136
rect 494244 700188 494296 700194
rect 494244 700130 494296 700136
rect 494796 700188 494848 700194
rect 494796 700130 494848 700136
rect 477880 698170 477908 700130
rect 494256 698170 494284 700130
rect 510632 699802 510660 703582
rect 510816 703474 510844 703582
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 511000 703474 511028 703520
rect 510816 703446 511028 703474
rect 527192 699802 527220 703520
rect 543476 702434 543504 703520
rect 559668 702434 559696 703520
rect 510540 699774 510660 699802
rect 526916 699774 527220 699802
rect 543200 702406 543504 702434
rect 559576 702406 559696 702434
rect 510540 698170 510568 699774
rect 526916 698170 526944 699774
rect 543200 698170 543228 702406
rect 559576 698170 559604 702406
rect 298020 698142 298092 698170
rect 216368 697959 216396 698142
rect 232744 697959 232772 698142
rect 249028 697959 249056 698142
rect 265404 697959 265432 698142
rect 281780 697959 281808 698142
rect 298064 697959 298092 698142
rect 314440 698142 314516 698170
rect 330724 698142 330800 698170
rect 347100 698142 347176 698170
rect 363476 698142 363552 698170
rect 379760 698142 379836 698170
rect 396136 698142 396212 698170
rect 412420 698142 412496 698170
rect 428796 698142 428872 698170
rect 445172 698142 445248 698170
rect 461456 698142 461532 698170
rect 477832 698142 477908 698170
rect 494208 698142 494284 698170
rect 510492 698142 510568 698170
rect 526868 698142 526944 698170
rect 543152 698142 543228 698170
rect 559528 698142 559604 698170
rect 575860 698170 575888 703520
rect 575860 698142 575932 698170
rect 314440 697959 314468 698142
rect 330724 697959 330752 698142
rect 347100 697959 347128 698142
rect 363476 697959 363504 698142
rect 379760 697959 379788 698142
rect 396136 697959 396164 698142
rect 412420 697959 412448 698142
rect 428796 697959 428824 698142
rect 445172 697959 445200 698142
rect 461456 697959 461484 698142
rect 477832 697959 477860 698142
rect 494208 697959 494236 698142
rect 510492 697959 510520 698142
rect 526868 697959 526896 698142
rect 543152 697959 543180 698142
rect 559528 697959 559556 698142
rect 575904 697959 575932 698142
rect 3514 697911 3570 697920
rect 3528 697377 3556 697911
rect 3514 697368 3570 697377
rect 3514 697303 3570 697312
rect 579526 684720 579582 684729
rect 579582 684678 579660 684706
rect 579526 684655 579582 684664
rect 579632 683913 579660 684678
rect 579618 683904 579674 683913
rect 579618 683839 579674 683848
rect 578330 644600 578386 644609
rect 578330 644535 578332 644544
rect 578384 644535 578386 644544
rect 580908 644564 580960 644570
rect 578332 644506 578384 644512
rect 580908 644506 580960 644512
rect 580920 644065 580948 644506
rect 580906 644056 580962 644065
rect 580906 643991 580962 644000
rect 3422 436656 3478 436665
rect 3422 436591 3478 436600
rect 3436 436051 3464 436591
rect 3422 436042 3478 436051
rect 3422 435977 3478 435986
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422997 3464 423535
rect 3422 422988 3478 422997
rect 3422 422923 3478 422932
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3436 409943 3464 410479
rect 3422 409934 3478 409943
rect 3422 409869 3478 409878
rect 3422 397488 3478 397497
rect 3422 397423 3478 397432
rect 3436 396889 3464 397423
rect 3422 396880 3478 396889
rect 3422 396815 3478 396824
rect 3422 384432 3478 384441
rect 3422 384367 3478 384376
rect 3436 383713 3464 384367
rect 3422 383704 3478 383713
rect 3422 383639 3478 383648
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 370659 3464 371311
rect 3422 370650 3478 370659
rect 3422 370585 3478 370594
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3436 357605 3464 358391
rect 3422 357596 3478 357605
rect 3422 357531 3478 357540
rect 579526 351928 579582 351937
rect 579526 351863 579582 351872
rect 579540 351121 579568 351863
rect 579526 351112 579582 351121
rect 579526 351047 579582 351056
rect 3422 345400 3478 345409
rect 3422 345335 3478 345344
rect 3436 344429 3464 345335
rect 3422 344420 3478 344429
rect 3422 344355 3478 344364
rect 579618 338600 579674 338609
rect 579618 338535 579674 338544
rect 579526 337920 579582 337929
rect 579632 337906 579660 338535
rect 579582 337878 579660 337906
rect 579526 337855 579582 337864
rect 3422 332344 3478 332353
rect 3422 332279 3478 332288
rect 3436 331375 3464 332279
rect 3422 331366 3478 331375
rect 3422 331301 3478 331310
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324465 580212 325207
rect 580170 324456 580226 324465
rect 580170 324391 580226 324400
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318321 3464 319223
rect 3422 318312 3478 318321
rect 3422 318247 3478 318256
rect 579618 312080 579674 312089
rect 579618 312015 579674 312024
rect 579526 311128 579582 311137
rect 579632 311114 579660 312015
rect 579582 311086 579660 311114
rect 579526 311063 579582 311072
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3436 305145 3464 306167
rect 3422 305136 3478 305145
rect 3422 305071 3478 305080
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 579526 297800 579582 297809
rect 579632 297786 579660 298687
rect 579582 297758 579660 297786
rect 579526 297735 579582 297744
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292091 3464 293111
rect 3422 292082 3478 292091
rect 3422 292017 3478 292026
rect 580170 285424 580226 285433
rect 580170 285359 580226 285368
rect 580184 284481 580212 285359
rect 580170 284472 580226 284481
rect 580170 284407 580226 284416
rect 3422 280120 3478 280129
rect 3422 280055 3478 280064
rect 3436 279037 3464 280055
rect 3422 279028 3478 279037
rect 3422 278963 3478 278972
rect 579618 272232 579674 272241
rect 579618 272167 579674 272176
rect 579526 271144 579582 271153
rect 579632 271130 579660 272167
rect 579582 271102 579660 271130
rect 579526 271079 579582 271088
rect 3422 267200 3478 267209
rect 3422 267135 3478 267144
rect 3436 265983 3464 267135
rect 3422 265974 3478 265983
rect 3422 265909 3478 265918
rect 580906 258904 580962 258913
rect 580906 258839 580962 258848
rect 580920 257854 580948 258839
rect 578884 257848 578936 257854
rect 578884 257790 578936 257796
rect 580908 257848 580960 257854
rect 580908 257790 580960 257796
rect 578896 257689 578924 257790
rect 578882 257680 578938 257689
rect 578882 257615 578938 257624
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 252807 3464 254079
rect 3422 252798 3478 252807
rect 3422 252733 3478 252742
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244497 580212 245511
rect 580170 244488 580226 244497
rect 580170 244423 580226 244432
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3436 239753 3464 241023
rect 3422 239744 3478 239753
rect 3422 239679 3478 239688
rect 579618 232384 579674 232393
rect 579618 232319 579674 232328
rect 579526 231160 579582 231169
rect 579632 231146 579660 232319
rect 579582 231118 579660 231146
rect 579526 231095 579582 231104
rect 3422 228032 3478 228041
rect 3422 227967 3478 227976
rect 3436 226699 3464 227967
rect 3422 226690 3478 226699
rect 3422 226625 3478 226634
rect 579618 219056 579674 219065
rect 579618 218991 579674 219000
rect 579526 217696 579582 217705
rect 579632 217682 579660 218991
rect 579582 217654 579660 217682
rect 579526 217631 579582 217640
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3436 213523 3464 214911
rect 3422 213514 3478 213523
rect 3422 213449 3478 213458
rect 579618 205728 579674 205737
rect 579618 205663 579674 205672
rect 579526 204368 579582 204377
rect 579632 204354 579660 205663
rect 579582 204326 579660 204354
rect 579526 204303 579582 204312
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3436 200469 3464 201855
rect 3422 200460 3478 200469
rect 3422 200395 3478 200404
rect 579618 192536 579674 192545
rect 579618 192471 579674 192480
rect 579526 191040 579582 191049
rect 579632 191026 579660 192471
rect 579582 190998 579660 191026
rect 579526 190975 579582 190984
rect 3606 188864 3662 188873
rect 3606 188799 3662 188808
rect 3620 187415 3648 188799
rect 3606 187406 3662 187415
rect 3606 187341 3662 187350
rect 579618 179208 579674 179217
rect 579618 179143 579674 179152
rect 579526 177712 579582 177721
rect 579632 177698 579660 179143
rect 579582 177670 579660 177698
rect 579526 177647 579582 177656
rect 3422 175944 3478 175953
rect 3422 175879 3478 175888
rect 3436 174239 3464 175879
rect 3422 174230 3478 174239
rect 3422 174165 3478 174174
rect 579618 165880 579674 165889
rect 579618 165815 579674 165824
rect 579526 164384 579582 164393
rect 579632 164370 579660 165815
rect 579582 164342 579660 164370
rect 579526 164319 579582 164328
rect 2134 162888 2190 162897
rect 2134 162823 2190 162832
rect 2148 161129 2176 162823
rect 2134 161120 2190 161129
rect 2134 161055 2190 161064
rect 580906 152688 580962 152697
rect 580906 152623 580962 152632
rect 580920 151502 580948 152623
rect 578516 151496 578568 151502
rect 578516 151438 578568 151444
rect 580908 151496 580960 151502
rect 580908 151438 580960 151444
rect 578528 151065 578556 151438
rect 578514 151056 578570 151065
rect 578514 150991 578570 151000
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3436 148131 3464 149767
rect 3422 148122 3478 148131
rect 3422 148057 3478 148066
rect 579618 139360 579674 139369
rect 579618 139295 579674 139304
rect 579526 137592 579582 137601
rect 579632 137578 579660 139295
rect 579582 137550 579660 137578
rect 579526 137527 579582 137536
rect 2134 136776 2190 136785
rect 2134 136711 2190 136720
rect 2148 135017 2176 136711
rect 2134 135008 2190 135017
rect 2134 134943 2190 134952
rect 579618 126032 579674 126041
rect 579618 125967 579674 125976
rect 579526 124400 579582 124409
rect 579632 124386 579660 125967
rect 579582 124358 579660 124386
rect 579526 124335 579582 124344
rect 3422 123720 3478 123729
rect 3422 123655 3478 123664
rect 3436 121901 3464 123655
rect 3422 121892 3478 121901
rect 3422 121827 3478 121836
rect 579618 112840 579674 112849
rect 579618 112775 579674 112784
rect 579526 110936 579582 110945
rect 579632 110922 579660 112775
rect 579582 110894 579660 110922
rect 579526 110871 579582 110880
rect 2134 110664 2190 110673
rect 2134 110599 2190 110608
rect 2148 108905 2176 110599
rect 2134 108896 2190 108905
rect 2134 108831 2190 108840
rect 579618 99512 579674 99521
rect 579618 99447 579674 99456
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 579526 97608 579582 97617
rect 579632 97594 579660 99447
rect 579582 97566 579660 97594
rect 579526 97543 579582 97552
rect 3436 95793 3464 97543
rect 3422 95784 3478 95793
rect 3422 95719 3478 95728
rect 579618 86184 579674 86193
rect 579618 86119 579674 86128
rect 2134 84688 2190 84697
rect 2134 84623 2190 84632
rect 2148 82657 2176 84623
rect 579526 84280 579582 84289
rect 579632 84266 579660 86119
rect 579582 84238 579660 84266
rect 579526 84215 579582 84224
rect 2134 82648 2190 82657
rect 2134 82583 2190 82592
rect 579618 72992 579674 73001
rect 579618 72927 579674 72936
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3436 69563 3464 71567
rect 579526 70952 579582 70961
rect 579632 70938 579660 72927
rect 579582 70910 579660 70938
rect 579526 70887 579582 70896
rect 3422 69554 3478 69563
rect 3422 69489 3478 69498
rect 579618 59664 579674 59673
rect 579618 59599 579674 59608
rect 2134 58576 2190 58585
rect 2134 58511 2190 58520
rect 2148 56545 2176 58511
rect 579526 57624 579582 57633
rect 579632 57610 579660 59599
rect 579582 57582 579660 57610
rect 579526 57559 579582 57568
rect 2134 56536 2190 56545
rect 2134 56471 2190 56480
rect 579986 46336 580042 46345
rect 579986 46271 580042 46280
rect 3422 45520 3478 45529
rect 3422 45455 3478 45464
rect 3436 43333 3464 45455
rect 580000 45014 580028 46271
rect 578332 45008 578384 45014
rect 578332 44950 578384 44956
rect 579988 45008 580040 45014
rect 579988 44950 580040 44956
rect 578344 44305 578372 44950
rect 578330 44296 578386 44305
rect 578330 44231 578386 44240
rect 3422 43324 3478 43333
rect 3422 43259 3478 43268
rect 579618 33144 579674 33153
rect 579618 33079 579674 33088
rect 2134 32464 2190 32473
rect 2134 32399 2190 32408
rect 2148 30297 2176 32399
rect 579526 30968 579582 30977
rect 579632 30954 579660 33079
rect 579582 30926 579660 30954
rect 579526 30903 579582 30912
rect 2134 30288 2190 30297
rect 2134 30223 2190 30232
rect 579618 19816 579674 19825
rect 579618 19751 579674 19760
rect 2042 19408 2098 19417
rect 2042 19343 2098 19352
rect 2056 17241 2084 19343
rect 579526 17640 579582 17649
rect 579632 17626 579660 19751
rect 579582 17598 579660 17626
rect 579526 17575 579582 17584
rect 2042 17232 2098 17241
rect 2042 17167 2098 17176
rect 579618 6624 579674 6633
rect 579618 6559 579674 6568
rect 2778 6488 2834 6497
rect 2778 6423 2834 6432
rect 2792 4185 2820 6423
rect 2778 4176 2834 4185
rect 2778 4111 2834 4120
rect 579526 4176 579582 4185
rect 579632 4162 579660 6559
rect 579582 4134 579660 4162
rect 579526 4111 579582 4120
rect 1676 3868 1728 3874
rect 1676 3810 1728 3816
rect 572 3800 624 3806
rect 572 3742 624 3748
rect 584 480 612 3742
rect 1688 480 1716 3810
rect 4124 3806 4152 4012
rect 5228 3874 5256 4012
rect 5216 3868 5268 3874
rect 5216 3810 5268 3816
rect 4112 3800 4164 3806
rect 6424 3754 6452 4012
rect 7528 3754 7556 4012
rect 4112 3742 4164 3748
rect 6380 3726 6452 3754
rect 7484 3726 7556 3754
rect 7656 3800 7708 3806
rect 8724 3754 8752 4012
rect 9920 3754 9948 4012
rect 11024 3806 11052 4012
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 7656 3742 7708 3748
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 3240 1352 3292 1358
rect 3240 1294 3292 1300
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 354 2954 480
rect 3252 354 3280 1294
rect 4080 480 4108 2858
rect 6380 1358 6408 3726
rect 7484 2922 7512 3726
rect 7472 2916 7524 2922
rect 7472 2858 7524 2864
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 5632 1148 5684 1154
rect 5632 1090 5684 1096
rect 2842 326 3280 354
rect 2842 -960 2954 326
rect 4038 -960 4150 480
rect 5234 354 5346 480
rect 5644 354 5672 1090
rect 6472 480 6500 2790
rect 7668 480 7696 3742
rect 8680 3726 8752 3754
rect 9876 3726 9948 3754
rect 11012 3800 11064 3806
rect 11012 3742 11064 3748
rect 8680 1154 8708 3726
rect 9876 2854 9904 3726
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 8668 1148 8720 1154
rect 8668 1090 8720 1096
rect 8760 944 8812 950
rect 8760 886 8812 892
rect 8772 480 8800 886
rect 9968 480 9996 2790
rect 11164 480 11192 3878
rect 12220 3754 12248 4012
rect 12176 3726 12248 3754
rect 12348 3800 12400 3806
rect 13324 3754 13352 4012
rect 14520 3942 14548 4012
rect 14508 3936 14560 3942
rect 14508 3878 14560 3884
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 13544 3868 13596 3874
rect 13544 3810 13596 3816
rect 12348 3742 12400 3748
rect 12176 950 12204 3726
rect 12164 944 12216 950
rect 12164 886 12216 892
rect 12360 480 12388 3742
rect 13280 3726 13352 3754
rect 13280 2854 13308 3726
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13556 480 13584 3810
rect 14752 480 14780 3878
rect 15716 3806 15744 4012
rect 16820 3874 16848 4012
rect 18016 3942 18044 4012
rect 18004 3936 18056 3942
rect 18004 3878 18056 3884
rect 16808 3868 16860 3874
rect 16808 3810 16860 3816
rect 19120 3806 19148 4012
rect 19432 3868 19484 3874
rect 19432 3810 19484 3816
rect 15704 3800 15756 3806
rect 15704 3742 15756 3748
rect 15936 3800 15988 3806
rect 15936 3742 15988 3748
rect 19108 3800 19160 3806
rect 19108 3742 19160 3748
rect 15948 480 15976 3742
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17052 480 17080 2790
rect 18248 480 18276 2858
rect 19444 480 19472 3810
rect 20316 3754 20344 4012
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20272 3726 20344 3754
rect 20272 2854 20300 3726
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 20640 480 20668 3878
rect 21512 3754 21540 4012
rect 22616 3874 22644 4012
rect 23812 3942 23840 4012
rect 23800 3936 23852 3942
rect 23800 3878 23852 3884
rect 24216 3936 24268 3942
rect 24216 3878 24268 3884
rect 22604 3868 22656 3874
rect 22604 3810 22656 3816
rect 23020 3868 23072 3874
rect 23020 3810 23072 3816
rect 21468 3726 21540 3754
rect 21824 3800 21876 3806
rect 21824 3742 21876 3748
rect 21468 2922 21496 3726
rect 21456 2916 21508 2922
rect 21456 2858 21508 2864
rect 21836 480 21864 3742
rect 23032 480 23060 3810
rect 24228 480 24256 3878
rect 24916 3806 24944 4012
rect 26112 3874 26140 4012
rect 27308 3942 27336 4012
rect 27296 3936 27348 3942
rect 27296 3878 27348 3884
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 26100 3868 26152 3874
rect 26100 3810 26152 3816
rect 26516 3868 26568 3874
rect 26516 3810 26568 3816
rect 24904 3800 24956 3806
rect 24904 3742 24956 3748
rect 25320 3800 25372 3806
rect 25320 3742 25372 3748
rect 25332 480 25360 3742
rect 26528 480 26556 3810
rect 27724 480 27752 3878
rect 28412 3806 28440 4012
rect 29608 3874 29636 4012
rect 30712 3942 30740 4012
rect 30700 3936 30752 3942
rect 30700 3878 30752 3884
rect 29596 3868 29648 3874
rect 29596 3810 29648 3816
rect 30104 3868 30156 3874
rect 30104 3810 30156 3816
rect 28400 3800 28452 3806
rect 28400 3742 28452 3748
rect 28908 2848 28960 2854
rect 28908 2790 28960 2796
rect 28920 480 28948 2790
rect 30116 480 30144 3810
rect 31300 3800 31352 3806
rect 31908 3754 31936 4012
rect 32404 3936 32456 3942
rect 32404 3878 32456 3884
rect 31300 3742 31352 3748
rect 31312 480 31340 3742
rect 31864 3726 31936 3754
rect 31864 2854 31892 3726
rect 31852 2848 31904 2854
rect 31852 2790 31904 2796
rect 32416 480 32444 3878
rect 33104 3874 33132 4012
rect 33092 3868 33144 3874
rect 33092 3810 33144 3816
rect 33600 3868 33652 3874
rect 33600 3810 33652 3816
rect 33612 480 33640 3810
rect 34208 3806 34236 4012
rect 35404 3942 35432 4012
rect 35392 3936 35444 3942
rect 35392 3878 35444 3884
rect 36600 3874 36628 4012
rect 36588 3868 36640 3874
rect 36588 3810 36640 3816
rect 37188 3868 37240 3874
rect 37188 3810 37240 3816
rect 34196 3800 34248 3806
rect 34196 3742 34248 3748
rect 34796 3800 34848 3806
rect 34796 3742 34848 3748
rect 34808 480 34836 3742
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 36004 480 36032 2790
rect 37200 480 37228 3810
rect 37704 3806 37732 4012
rect 38384 3936 38436 3942
rect 38384 3878 38436 3884
rect 37692 3800 37744 3806
rect 37692 3742 37744 3748
rect 38396 480 38424 3878
rect 38900 3754 38928 4012
rect 40004 3874 40032 4012
rect 41200 3942 41228 4012
rect 41188 3936 41240 3942
rect 41188 3878 41240 3884
rect 39992 3868 40044 3874
rect 39992 3810 40044 3816
rect 41880 3868 41932 3874
rect 41880 3810 41932 3816
rect 38856 3726 38928 3754
rect 40684 3800 40736 3806
rect 40684 3742 40736 3748
rect 38856 2854 38884 3726
rect 38844 2848 38896 2854
rect 38844 2790 38896 2796
rect 39580 2848 39632 2854
rect 39580 2790 39632 2796
rect 39592 480 39620 2790
rect 40696 480 40724 3742
rect 41892 480 41920 3810
rect 42396 3754 42424 4012
rect 43076 3936 43128 3942
rect 43076 3878 43128 3884
rect 42352 3726 42424 3754
rect 42352 2854 42380 3726
rect 42340 2848 42392 2854
rect 42340 2790 42392 2796
rect 43088 480 43116 3878
rect 43500 3806 43528 4012
rect 44696 3874 44724 4012
rect 45800 3942 45828 4012
rect 45788 3936 45840 3942
rect 45788 3878 45840 3884
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 44684 3868 44736 3874
rect 44684 3810 44736 3816
rect 45468 3868 45520 3874
rect 45468 3810 45520 3816
rect 43488 3800 43540 3806
rect 43488 3742 43540 3748
rect 44272 3800 44324 3806
rect 44272 3742 44324 3748
rect 44284 480 44312 3742
rect 45480 480 45508 3810
rect 46676 480 46704 3878
rect 46996 3806 47024 4012
rect 48192 3874 48220 4012
rect 49296 3942 49324 4012
rect 49284 3936 49336 3942
rect 49284 3878 49336 3884
rect 50160 3936 50212 3942
rect 50160 3878 50212 3884
rect 48180 3868 48232 3874
rect 48180 3810 48232 3816
rect 48964 3868 49016 3874
rect 48964 3810 49016 3816
rect 46984 3800 47036 3806
rect 46984 3742 47036 3748
rect 47860 3800 47912 3806
rect 47860 3742 47912 3748
rect 47872 480 47900 3742
rect 48976 480 49004 3810
rect 50172 480 50200 3878
rect 50492 3806 50520 4012
rect 51596 3874 51624 4012
rect 52792 3942 52820 4012
rect 52780 3936 52832 3942
rect 52780 3878 52832 3884
rect 51584 3868 51636 3874
rect 51584 3810 51636 3816
rect 53748 3868 53800 3874
rect 53748 3810 53800 3816
rect 50480 3800 50532 3806
rect 50480 3742 50532 3748
rect 51356 3800 51408 3806
rect 51356 3742 51408 3748
rect 51368 480 51396 3742
rect 52552 740 52604 746
rect 52552 682 52604 688
rect 52564 480 52592 682
rect 53760 480 53788 3810
rect 53988 3806 54016 4012
rect 53976 3800 54028 3806
rect 53976 3742 54028 3748
rect 54944 3800 54996 3806
rect 55092 3754 55120 4012
rect 56048 3936 56100 3942
rect 56048 3878 56100 3884
rect 54944 3742 54996 3748
rect 54956 480 54984 3742
rect 55048 3726 55120 3754
rect 55048 746 55076 3726
rect 55036 740 55088 746
rect 55036 682 55088 688
rect 56060 480 56088 3878
rect 56288 3874 56316 4012
rect 56276 3868 56328 3874
rect 56276 3810 56328 3816
rect 57244 3868 57296 3874
rect 57244 3810 57296 3816
rect 57256 480 57284 3810
rect 57392 3806 57420 4012
rect 58588 3942 58616 4012
rect 58576 3936 58628 3942
rect 58576 3878 58628 3884
rect 59784 3874 59812 4012
rect 59772 3868 59824 3874
rect 59772 3810 59824 3816
rect 60888 3806 60916 4012
rect 62084 3890 62112 4012
rect 61948 3862 62112 3890
rect 57380 3800 57432 3806
rect 57380 3742 57432 3748
rect 58440 3800 58492 3806
rect 58440 3742 58492 3748
rect 60876 3800 60928 3806
rect 60876 3742 60928 3748
rect 58452 480 58480 3742
rect 60832 1352 60884 1358
rect 60832 1294 60884 1300
rect 59636 740 59688 746
rect 59636 682 59688 688
rect 59648 480 59676 682
rect 60844 480 60872 1294
rect 61948 746 61976 3862
rect 63280 3754 63308 4012
rect 64384 3890 64412 4012
rect 64384 3862 64460 3890
rect 64328 3800 64380 3806
rect 63280 3726 63356 3754
rect 64328 3742 64380 3748
rect 63224 3052 63276 3058
rect 63224 2994 63276 3000
rect 62028 2848 62080 2854
rect 62028 2790 62080 2796
rect 61936 740 61988 746
rect 61936 682 61988 688
rect 62040 480 62068 2790
rect 63236 480 63264 2994
rect 63328 1358 63356 3726
rect 63316 1352 63368 1358
rect 63316 1294 63368 1300
rect 64340 480 64368 3742
rect 64432 2854 64460 3862
rect 65580 3754 65608 4012
rect 66684 3806 66712 4012
rect 65536 3726 65608 3754
rect 66672 3800 66724 3806
rect 66672 3742 66724 3748
rect 67088 3800 67140 3806
rect 67880 3754 67908 4012
rect 69076 3806 69104 4012
rect 67088 3742 67140 3748
rect 65536 3058 65564 3726
rect 65524 3052 65576 3058
rect 65524 2994 65576 3000
rect 64420 2848 64472 2854
rect 64420 2790 64472 2796
rect 65524 2848 65576 2854
rect 65524 2790 65576 2796
rect 65536 480 65564 2790
rect 5234 326 5672 354
rect 5234 -960 5346 326
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 218 66802 480
rect 67100 218 67128 3742
rect 67836 3726 67908 3754
rect 69064 3800 69116 3806
rect 70180 3754 70208 4012
rect 69064 3742 69116 3748
rect 70136 3726 70208 3754
rect 70308 3800 70360 3806
rect 71376 3754 71404 4012
rect 71504 3868 71556 3874
rect 71504 3810 71556 3816
rect 70308 3742 70360 3748
rect 67836 2854 67864 3726
rect 67824 2848 67876 2854
rect 67824 2790 67876 2796
rect 70136 1358 70164 3726
rect 67916 1352 67968 1358
rect 67916 1294 67968 1300
rect 70124 1352 70176 1358
rect 70124 1294 70176 1300
rect 67928 480 67956 1294
rect 69112 604 69164 610
rect 69112 546 69164 552
rect 69124 480 69152 546
rect 70320 480 70348 3742
rect 71332 3726 71404 3754
rect 71332 610 71360 3726
rect 71320 604 71372 610
rect 71320 546 71372 552
rect 71516 480 71544 3810
rect 72480 3806 72508 4012
rect 72608 3936 72660 3942
rect 72608 3878 72660 3884
rect 72468 3800 72520 3806
rect 72468 3742 72520 3748
rect 72620 480 72648 3878
rect 73676 3874 73704 4012
rect 74872 3942 74900 4012
rect 74860 3936 74912 3942
rect 74860 3878 74912 3884
rect 73664 3868 73716 3874
rect 73664 3810 73716 3816
rect 75976 3806 76004 4012
rect 73804 3800 73856 3806
rect 73804 3742 73856 3748
rect 75964 3800 76016 3806
rect 77172 3754 77200 4012
rect 78276 3754 78304 4012
rect 78588 3868 78640 3874
rect 78588 3810 78640 3816
rect 75964 3742 76016 3748
rect 73816 480 73844 3742
rect 77128 3726 77200 3754
rect 78232 3726 78304 3754
rect 76196 1352 76248 1358
rect 76196 1294 76248 1300
rect 75000 1284 75052 1290
rect 75000 1226 75052 1232
rect 75012 480 75040 1226
rect 76208 480 76236 1294
rect 77128 1290 77156 3726
rect 78232 1358 78260 3726
rect 78220 1352 78272 1358
rect 78220 1294 78272 1300
rect 77116 1284 77168 1290
rect 77116 1226 77168 1232
rect 77392 1284 77444 1290
rect 77392 1226 77444 1232
rect 77404 480 77432 1226
rect 78600 480 78628 3810
rect 79472 3754 79500 4012
rect 80668 3874 80696 4012
rect 80656 3868 80708 3874
rect 80656 3810 80708 3816
rect 80888 3868 80940 3874
rect 80888 3810 80940 3816
rect 79428 3726 79500 3754
rect 79692 3800 79744 3806
rect 79692 3742 79744 3748
rect 79428 1290 79456 3726
rect 79416 1284 79468 1290
rect 79416 1226 79468 1232
rect 79704 480 79732 3742
rect 80900 480 80928 3810
rect 81772 3806 81800 4012
rect 82968 3874 82996 4012
rect 82956 3868 83008 3874
rect 82956 3810 83008 3816
rect 81760 3800 81812 3806
rect 84072 3754 84100 4012
rect 85268 3754 85296 4012
rect 86464 3754 86492 4012
rect 81760 3742 81812 3748
rect 84028 3726 84100 3754
rect 85224 3726 85296 3754
rect 86420 3726 86492 3754
rect 86868 3800 86920 3806
rect 87568 3754 87596 4012
rect 87972 3868 88024 3874
rect 87972 3810 88024 3816
rect 86868 3742 86920 3748
rect 83280 1352 83332 1358
rect 83280 1294 83332 1300
rect 82084 1284 82136 1290
rect 82084 1226 82136 1232
rect 82096 480 82124 1226
rect 83292 480 83320 1294
rect 84028 1290 84056 3726
rect 85224 1358 85252 3726
rect 85212 1352 85264 1358
rect 85212 1294 85264 1300
rect 85672 1352 85724 1358
rect 85672 1294 85724 1300
rect 84016 1284 84068 1290
rect 84016 1226 84068 1232
rect 84476 1284 84528 1290
rect 84476 1226 84528 1232
rect 84488 480 84516 1226
rect 85684 480 85712 1294
rect 86420 1290 86448 3726
rect 86408 1284 86460 1290
rect 86408 1226 86460 1232
rect 86880 480 86908 3742
rect 87524 3726 87596 3754
rect 87524 1358 87552 3726
rect 87512 1352 87564 1358
rect 87512 1294 87564 1300
rect 87984 480 88012 3810
rect 88764 3806 88792 4012
rect 89960 3874 89988 4012
rect 89948 3868 90000 3874
rect 89948 3810 90000 3816
rect 88752 3800 88804 3806
rect 91064 3754 91092 4012
rect 92260 3754 92288 4012
rect 93364 3754 93392 4012
rect 94560 3754 94588 4012
rect 88752 3742 88804 3748
rect 91020 3726 91092 3754
rect 92216 3726 92288 3754
rect 93320 3726 93392 3754
rect 94516 3726 94588 3754
rect 95148 3800 95200 3806
rect 95756 3754 95784 4012
rect 96252 3868 96304 3874
rect 96252 3810 96304 3816
rect 95148 3742 95200 3748
rect 91020 1358 91048 3726
rect 89168 1352 89220 1358
rect 89168 1294 89220 1300
rect 91008 1352 91060 1358
rect 91008 1294 91060 1300
rect 91560 1352 91612 1358
rect 91560 1294 91612 1300
rect 89180 480 89208 1294
rect 90364 1284 90416 1290
rect 90364 1226 90416 1232
rect 90376 480 90404 1226
rect 91572 480 91600 1294
rect 92216 1290 92244 3726
rect 93320 1358 93348 3726
rect 93308 1352 93360 1358
rect 93308 1294 93360 1300
rect 93952 1352 94004 1358
rect 93952 1294 94004 1300
rect 92204 1284 92256 1290
rect 92204 1226 92256 1232
rect 92756 1284 92808 1290
rect 92756 1226 92808 1232
rect 92768 480 92796 1226
rect 93964 480 93992 1294
rect 94516 1290 94544 3726
rect 94504 1284 94556 1290
rect 94504 1226 94556 1232
rect 95160 480 95188 3742
rect 95712 3726 95784 3754
rect 95712 1358 95740 3726
rect 95700 1352 95752 1358
rect 95700 1294 95752 1300
rect 96264 480 96292 3810
rect 96860 3806 96888 4012
rect 98056 3874 98084 4012
rect 98044 3868 98096 3874
rect 98044 3810 98096 3816
rect 96848 3800 96900 3806
rect 99160 3754 99188 4012
rect 100356 3754 100384 4012
rect 101552 3754 101580 4012
rect 102656 3754 102684 4012
rect 96848 3742 96900 3748
rect 99116 3726 99188 3754
rect 100312 3726 100384 3754
rect 101508 3726 101580 3754
rect 102612 3726 102684 3754
rect 103336 3800 103388 3806
rect 103852 3754 103880 4012
rect 104956 3806 104984 4012
rect 103336 3742 103388 3748
rect 99116 1358 99144 3726
rect 97448 1352 97500 1358
rect 97448 1294 97500 1300
rect 99104 1352 99156 1358
rect 99104 1294 99156 1300
rect 97460 480 97488 1294
rect 100312 1290 100340 3726
rect 101036 1352 101088 1358
rect 101036 1294 101088 1300
rect 98644 1284 98696 1290
rect 98644 1226 98696 1232
rect 100300 1284 100352 1290
rect 100300 1226 100352 1232
rect 98656 480 98684 1226
rect 99840 1216 99892 1222
rect 99840 1158 99892 1164
rect 99852 480 99880 1158
rect 101048 480 101076 1294
rect 101508 1222 101536 3726
rect 102612 1358 102640 3726
rect 102600 1352 102652 1358
rect 102600 1294 102652 1300
rect 102232 1284 102284 1290
rect 102232 1226 102284 1232
rect 101496 1216 101548 1222
rect 101496 1158 101548 1164
rect 102244 480 102272 1226
rect 103348 480 103376 3742
rect 103808 3726 103880 3754
rect 104944 3800 104996 3806
rect 106152 3754 106180 4012
rect 107348 3754 107376 4012
rect 108452 3754 108480 4012
rect 109648 3754 109676 4012
rect 110752 3754 110780 4012
rect 111948 3754 111976 4012
rect 113144 3754 113172 4012
rect 114248 3754 114276 4012
rect 115444 3754 115472 4012
rect 116640 3754 116668 4012
rect 117744 3754 117772 4012
rect 118940 3754 118968 4012
rect 120044 3754 120072 4012
rect 121240 3754 121268 4012
rect 122436 3754 122464 4012
rect 123540 3754 123568 4012
rect 104944 3742 104996 3748
rect 106108 3726 106180 3754
rect 107304 3726 107376 3754
rect 108408 3726 108480 3754
rect 109604 3726 109676 3754
rect 110708 3726 110780 3754
rect 111904 3726 111976 3754
rect 113100 3726 113172 3754
rect 114204 3726 114276 3754
rect 115400 3726 115472 3754
rect 116596 3726 116668 3754
rect 117700 3726 117772 3754
rect 118896 3726 118968 3754
rect 119264 3726 120072 3754
rect 121196 3726 121268 3754
rect 122392 3726 122464 3754
rect 123496 3726 123568 3754
rect 124736 3754 124764 4012
rect 125840 3754 125868 4012
rect 127036 3754 127064 4012
rect 128232 3754 128260 4012
rect 129336 3754 129364 4012
rect 130532 3754 130560 4012
rect 131636 3754 131664 4012
rect 132832 3754 132860 4012
rect 134028 3754 134056 4012
rect 135132 3754 135160 4012
rect 136328 3754 136356 4012
rect 137432 3754 137460 4012
rect 138628 3754 138656 4012
rect 139824 3754 139852 4012
rect 140928 3754 140956 4012
rect 142124 3754 142152 4012
rect 143320 3754 143348 4012
rect 144424 3754 144452 4012
rect 145620 3754 145648 4012
rect 146724 3754 146752 4012
rect 147920 3754 147948 4012
rect 149116 3754 149144 4012
rect 150220 3754 150248 4012
rect 151416 3754 151444 4012
rect 152520 3754 152548 4012
rect 153716 3754 153744 4012
rect 154912 3754 154940 4012
rect 156016 3754 156044 4012
rect 157212 3754 157240 4012
rect 158316 3754 158344 4012
rect 159512 3754 159540 4012
rect 160708 3754 160736 4012
rect 161812 3754 161840 4012
rect 163008 3754 163036 4012
rect 164112 3754 164140 4012
rect 165308 3754 165336 4012
rect 166504 3754 166532 4012
rect 167608 3754 167636 4012
rect 168804 3754 168832 4012
rect 170000 3754 170028 4012
rect 171104 3754 171132 4012
rect 172300 3754 172328 4012
rect 173404 3754 173432 4012
rect 174600 3754 174628 4012
rect 175796 3754 175824 4012
rect 176900 3754 176928 4012
rect 178096 3754 178124 4012
rect 179200 3754 179228 4012
rect 124736 3726 124812 3754
rect 103808 1290 103836 3726
rect 106108 1358 106136 3726
rect 104532 1352 104584 1358
rect 104532 1294 104584 1300
rect 106096 1352 106148 1358
rect 106096 1294 106148 1300
rect 106924 1352 106976 1358
rect 106924 1294 106976 1300
rect 103796 1284 103848 1290
rect 103796 1226 103848 1232
rect 104544 480 104572 1294
rect 105728 740 105780 746
rect 105728 682 105780 688
rect 105740 480 105768 682
rect 106936 480 106964 1294
rect 107304 746 107332 3726
rect 108408 1358 108436 3726
rect 108396 1352 108448 1358
rect 108396 1294 108448 1300
rect 109316 1352 109368 1358
rect 109316 1294 109368 1300
rect 108120 1284 108172 1290
rect 108120 1226 108172 1232
rect 107292 740 107344 746
rect 107292 682 107344 688
rect 108132 480 108160 1226
rect 109328 480 109356 1294
rect 109604 1290 109632 3726
rect 110708 1358 110736 3726
rect 110696 1352 110748 1358
rect 110696 1294 110748 1300
rect 111904 1290 111932 3726
rect 112812 1352 112864 1358
rect 112812 1294 112864 1300
rect 109592 1284 109644 1290
rect 109592 1226 109644 1232
rect 110512 1284 110564 1290
rect 110512 1226 110564 1232
rect 111892 1284 111944 1290
rect 111892 1226 111944 1232
rect 110524 480 110552 1226
rect 111616 1148 111668 1154
rect 111616 1090 111668 1096
rect 111628 480 111656 1090
rect 112824 480 112852 1294
rect 113100 1154 113128 3726
rect 114204 1358 114232 3726
rect 114192 1352 114244 1358
rect 114192 1294 114244 1300
rect 115204 1284 115256 1290
rect 115204 1226 115256 1232
rect 114008 1216 114060 1222
rect 114008 1158 114060 1164
rect 113088 1148 113140 1154
rect 113088 1090 113140 1096
rect 114020 480 114048 1158
rect 115216 480 115244 1226
rect 115400 1222 115428 3726
rect 116400 1352 116452 1358
rect 116400 1294 116452 1300
rect 115388 1216 115440 1222
rect 115388 1158 115440 1164
rect 116412 480 116440 1294
rect 116596 1290 116624 3726
rect 117700 1358 117728 3726
rect 117688 1352 117740 1358
rect 117688 1294 117740 1300
rect 118896 1290 118924 3726
rect 116584 1284 116636 1290
rect 116584 1226 116636 1232
rect 117596 1284 117648 1290
rect 117596 1226 117648 1232
rect 118884 1284 118936 1290
rect 118884 1226 118936 1232
rect 117608 480 117636 1226
rect 66690 190 67128 218
rect 66690 -960 66802 190
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 354 118874 480
rect 119264 354 119292 3726
rect 121196 1358 121224 3726
rect 119896 1352 119948 1358
rect 119896 1294 119948 1300
rect 121184 1352 121236 1358
rect 121184 1294 121236 1300
rect 119908 480 119936 1294
rect 122288 1284 122340 1290
rect 122288 1226 122340 1232
rect 121092 944 121144 950
rect 121092 886 121144 892
rect 121104 480 121132 886
rect 122300 480 122328 1226
rect 122392 950 122420 3726
rect 123496 1290 123524 3726
rect 123484 1284 123536 1290
rect 123484 1226 123536 1232
rect 124680 1284 124732 1290
rect 124680 1226 124732 1232
rect 123484 1148 123536 1154
rect 123484 1090 123536 1096
rect 122380 944 122432 950
rect 122380 886 122432 892
rect 123496 480 123524 1090
rect 124692 480 124720 1226
rect 124784 1154 124812 3726
rect 125796 3726 125868 3754
rect 126992 3726 127064 3754
rect 127176 3726 128260 3754
rect 129292 3726 129364 3754
rect 130488 3726 130560 3754
rect 131592 3726 131664 3754
rect 132788 3726 132860 3754
rect 133984 3726 134056 3754
rect 134168 3726 135160 3754
rect 135272 3726 136356 3754
rect 137388 3726 137460 3754
rect 138584 3726 138656 3754
rect 139780 3726 139852 3754
rect 140884 3726 140956 3754
rect 141712 3726 142152 3754
rect 142448 3726 143348 3754
rect 143552 3726 144452 3754
rect 145576 3726 145648 3754
rect 146680 3726 146752 3754
rect 147600 3726 147948 3754
rect 149072 3726 149144 3754
rect 149992 3726 150248 3754
rect 151096 3726 151444 3754
rect 151832 3726 152548 3754
rect 153488 3726 153744 3754
rect 154868 3726 154940 3754
rect 155880 3726 156044 3754
rect 156616 3726 157240 3754
rect 158272 3726 158344 3754
rect 159376 3726 159540 3754
rect 160112 3726 160736 3754
rect 161584 3726 161840 3754
rect 162964 3726 163036 3754
rect 164068 3726 164140 3754
rect 164896 3726 165336 3754
rect 166460 3726 166532 3754
rect 167564 3726 167636 3754
rect 168392 3726 168832 3754
rect 169956 3726 170028 3754
rect 170784 3726 171132 3754
rect 172256 3726 172328 3754
rect 173176 3726 173432 3754
rect 174280 3726 174628 3754
rect 175752 3726 175824 3754
rect 176672 3726 176928 3754
rect 178052 3726 178124 3754
rect 179064 3726 179228 3754
rect 180396 3754 180424 4012
rect 181592 3754 181620 4012
rect 182696 3754 182724 4012
rect 180396 3726 180472 3754
rect 125796 1290 125824 3726
rect 126992 1358 127020 3726
rect 125876 1352 125928 1358
rect 125876 1294 125928 1300
rect 126980 1352 127032 1358
rect 126980 1294 127032 1300
rect 125784 1284 125836 1290
rect 125784 1226 125836 1232
rect 124772 1148 124824 1154
rect 124772 1090 124824 1096
rect 125888 480 125916 1294
rect 127176 1170 127204 3726
rect 129292 1290 129320 3726
rect 130488 1358 130516 3726
rect 131592 1358 131620 3726
rect 132788 1358 132816 3726
rect 133984 1358 134012 3726
rect 129372 1352 129424 1358
rect 129372 1294 129424 1300
rect 130476 1352 130528 1358
rect 130476 1294 130528 1300
rect 130568 1352 130620 1358
rect 130568 1294 130620 1300
rect 131580 1352 131632 1358
rect 131580 1294 131632 1300
rect 131764 1352 131816 1358
rect 131764 1294 131816 1300
rect 132776 1352 132828 1358
rect 132776 1294 132828 1300
rect 132960 1352 133012 1358
rect 132960 1294 133012 1300
rect 133972 1352 134024 1358
rect 133972 1294 134024 1300
rect 128176 1284 128228 1290
rect 128176 1226 128228 1232
rect 129280 1284 129332 1290
rect 129280 1226 129332 1232
rect 126992 1142 127204 1170
rect 126992 480 127020 1142
rect 128188 480 128216 1226
rect 129384 480 129412 1294
rect 130580 480 130608 1294
rect 131776 480 131804 1294
rect 132972 480 133000 1294
rect 134168 480 134196 3726
rect 135272 480 135300 3726
rect 137388 1290 137416 3726
rect 138584 1358 138612 3726
rect 137652 1352 137704 1358
rect 137652 1294 137704 1300
rect 138572 1352 138624 1358
rect 138572 1294 138624 1300
rect 136456 1284 136508 1290
rect 136456 1226 136508 1232
rect 137376 1284 137428 1290
rect 137376 1226 137428 1232
rect 136468 480 136496 1226
rect 137664 480 137692 1294
rect 139780 1290 139808 3726
rect 140884 1290 140912 3726
rect 138848 1284 138900 1290
rect 138848 1226 138900 1232
rect 139768 1284 139820 1290
rect 139768 1226 139820 1232
rect 140044 1284 140096 1290
rect 140044 1226 140096 1232
rect 140872 1284 140924 1290
rect 140872 1226 140924 1232
rect 138860 480 138888 1226
rect 140056 480 140084 1226
rect 118762 326 119292 354
rect 118762 -960 118874 326
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 354 141322 480
rect 141712 354 141740 3726
rect 142448 480 142476 3726
rect 143552 480 143580 3726
rect 145576 1358 145604 3726
rect 146680 1358 146708 3726
rect 144736 1352 144788 1358
rect 144736 1294 144788 1300
rect 145564 1352 145616 1358
rect 145564 1294 145616 1300
rect 145932 1352 145984 1358
rect 145932 1294 145984 1300
rect 146668 1352 146720 1358
rect 146668 1294 146720 1300
rect 144748 480 144776 1294
rect 145944 480 145972 1294
rect 141210 326 141740 354
rect 141210 -960 141322 326
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 354 147210 480
rect 147600 354 147628 3726
rect 149072 1358 149100 3726
rect 148324 1352 148376 1358
rect 148324 1294 148376 1300
rect 149060 1352 149112 1358
rect 149060 1294 149112 1300
rect 148336 480 148364 1294
rect 147098 326 147628 354
rect 147098 -960 147210 326
rect 148294 -960 148406 480
rect 149490 354 149602 480
rect 149992 354 150020 3726
rect 149490 326 150020 354
rect 150594 354 150706 480
rect 151096 354 151124 3726
rect 151832 480 151860 3726
rect 150594 326 151124 354
rect 149490 -960 149602 326
rect 150594 -960 150706 326
rect 151790 -960 151902 480
rect 152986 354 153098 480
rect 153488 354 153516 3726
rect 154868 1358 154896 3726
rect 154212 1352 154264 1358
rect 154212 1294 154264 1300
rect 154856 1352 154908 1358
rect 154856 1294 154908 1300
rect 154224 480 154252 1294
rect 152986 326 153516 354
rect 152986 -960 153098 326
rect 154182 -960 154294 480
rect 155378 354 155490 480
rect 155880 354 155908 3726
rect 156616 480 156644 3726
rect 155378 326 155908 354
rect 155378 -960 155490 326
rect 156574 -960 156686 480
rect 157770 354 157882 480
rect 158272 354 158300 3726
rect 157770 326 158300 354
rect 158874 354 158986 480
rect 159376 354 159404 3726
rect 160112 480 160140 3726
rect 158874 326 159404 354
rect 157770 -960 157882 326
rect 158874 -960 158986 326
rect 160070 -960 160182 480
rect 161266 354 161378 480
rect 161584 354 161612 3726
rect 162964 1358 162992 3726
rect 162492 1352 162544 1358
rect 162492 1294 162544 1300
rect 162952 1352 163004 1358
rect 162952 1294 163004 1300
rect 162504 480 162532 1294
rect 161266 326 161612 354
rect 161266 -960 161378 326
rect 162462 -960 162574 480
rect 163658 354 163770 480
rect 164068 354 164096 3726
rect 164896 480 164924 3726
rect 163658 326 164096 354
rect 163658 -960 163770 326
rect 164854 -960 164966 480
rect 166050 354 166162 480
rect 166460 354 166488 3726
rect 166050 326 166488 354
rect 167154 354 167266 480
rect 167564 354 167592 3726
rect 168392 480 168420 3726
rect 167154 326 167592 354
rect 166050 -960 166162 326
rect 167154 -960 167266 326
rect 168350 -960 168462 480
rect 169546 354 169658 480
rect 169956 354 169984 3726
rect 170784 480 170812 3726
rect 169546 326 169984 354
rect 169546 -960 169658 326
rect 170742 -960 170854 480
rect 171938 354 172050 480
rect 172256 354 172284 3726
rect 173176 480 173204 3726
rect 174280 480 174308 3726
rect 171938 326 172284 354
rect 171938 -960 172050 326
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 354 175546 480
rect 175752 354 175780 3726
rect 176672 480 176700 3726
rect 175434 326 175780 354
rect 175434 -960 175546 326
rect 176630 -960 176742 480
rect 177826 354 177938 480
rect 178052 354 178080 3726
rect 179064 480 179092 3726
rect 177826 326 178080 354
rect 177826 -960 177938 326
rect 179022 -960 179134 480
rect 180218 218 180330 480
rect 180444 218 180472 3726
rect 181456 3726 181620 3754
rect 182560 3726 182724 3754
rect 183892 3754 183920 4012
rect 184996 3754 185024 4012
rect 186192 3754 186220 4012
rect 187388 3754 187416 4012
rect 183892 3726 183968 3754
rect 181456 480 181484 3726
rect 182560 480 182588 3726
rect 180218 190 180472 218
rect 180218 -960 180330 190
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 218 183826 480
rect 183940 218 183968 3726
rect 184952 3726 185024 3754
rect 186148 3726 186220 3754
rect 187344 3726 187416 3754
rect 188492 3754 188520 4012
rect 189688 3754 189716 4012
rect 190792 3754 190820 4012
rect 191988 3754 192016 4012
rect 193184 3754 193212 4012
rect 194288 3754 194316 4012
rect 195484 3754 195512 4012
rect 188492 3726 188568 3754
rect 189688 3726 189764 3754
rect 190792 3726 190868 3754
rect 191988 3726 192064 3754
rect 193184 3726 193260 3754
rect 194288 3726 194456 3754
rect 184952 480 184980 3726
rect 186148 480 186176 3726
rect 187344 480 187372 3726
rect 188540 480 188568 3726
rect 189736 480 189764 3726
rect 190840 480 190868 3726
rect 192036 480 192064 3726
rect 193232 480 193260 3726
rect 194428 480 194456 3726
rect 195440 3726 195512 3754
rect 196680 3754 196708 4012
rect 197784 3754 197812 4012
rect 198980 3754 199008 4012
rect 196680 3726 196848 3754
rect 197784 3726 197952 3754
rect 183714 190 183968 218
rect 183714 -960 183826 190
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195440 218 195468 3726
rect 196820 480 196848 3726
rect 197924 480 197952 3726
rect 198936 3726 199008 3754
rect 200084 3754 200112 4012
rect 201280 3754 201308 4012
rect 202476 3754 202504 4012
rect 203580 3754 203608 4012
rect 204776 3754 204804 4012
rect 205880 3754 205908 4012
rect 207076 3754 207104 4012
rect 208272 3754 208300 4012
rect 209376 3754 209404 4012
rect 210572 3754 210600 4012
rect 211676 3754 211704 4012
rect 212872 3754 212900 4012
rect 214068 3754 214096 4012
rect 215172 3754 215200 4012
rect 216368 3806 216396 4012
rect 216356 3800 216408 3806
rect 200084 3726 200344 3754
rect 201280 3726 201356 3754
rect 202476 3726 202736 3754
rect 203580 3726 203656 3754
rect 204776 3726 205128 3754
rect 205880 3726 206232 3754
rect 207076 3726 207152 3754
rect 208272 3726 208624 3754
rect 209376 3726 209728 3754
rect 210572 3726 211016 3754
rect 211676 3726 211752 3754
rect 212872 3726 213408 3754
rect 214068 3726 214512 3754
rect 215172 3726 215248 3754
rect 216356 3742 216408 3748
rect 216864 3800 216916 3806
rect 216864 3742 216916 3748
rect 217472 3754 217500 4012
rect 218668 3754 218696 4012
rect 219864 3754 219892 4012
rect 220968 3754 220996 4012
rect 222164 3806 222192 4012
rect 222152 3800 222204 3806
rect 195582 218 195694 480
rect 195440 190 195694 218
rect 195582 -960 195694 190
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198936 218 198964 3726
rect 200316 480 200344 3726
rect 199078 218 199190 480
rect 198936 190 199190 218
rect 199078 -960 199190 190
rect 200274 -960 200386 480
rect 201328 354 201356 3726
rect 202708 480 202736 3726
rect 201470 354 201582 480
rect 201328 326 201582 354
rect 201470 -960 201582 326
rect 202666 -960 202778 480
rect 203628 354 203656 3726
rect 205100 480 205128 3726
rect 206204 480 206232 3726
rect 203862 354 203974 480
rect 203628 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207124 354 207152 3726
rect 208596 480 208624 3726
rect 209700 626 209728 3726
rect 209700 598 209774 626
rect 209746 480 209774 598
rect 210988 480 211016 3726
rect 207358 354 207470 480
rect 207124 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209746 326 209862 480
rect 209750 -960 209862 326
rect 210946 -960 211058 480
rect 211724 354 211752 3726
rect 213380 480 213408 3726
rect 214484 480 214512 3726
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215220 354 215248 3726
rect 216876 480 216904 3742
rect 217472 3726 217640 3754
rect 218668 3726 219296 3754
rect 219864 3726 220032 3754
rect 220968 3726 221136 3754
rect 222152 3742 222204 3748
rect 222752 3800 222804 3806
rect 222752 3742 222804 3748
rect 223360 3754 223388 4012
rect 224464 3806 224492 4012
rect 224452 3800 224504 3806
rect 215638 354 215750 480
rect 215220 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 217612 354 217640 3726
rect 219268 480 219296 3726
rect 218030 354 218142 480
rect 217612 326 218142 354
rect 218030 -960 218142 326
rect 219226 -960 219338 480
rect 220004 354 220032 3726
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 3726
rect 222764 480 222792 3742
rect 223360 3726 223528 3754
rect 224452 3742 224504 3748
rect 225144 3800 225196 3806
rect 225144 3742 225196 3748
rect 225660 3754 225688 4012
rect 226764 3754 226792 4012
rect 227960 3754 227988 4012
rect 229156 3754 229184 4012
rect 230260 3806 230288 4012
rect 231456 3806 231484 4012
rect 232560 3806 232588 4012
rect 233756 3806 233784 4012
rect 230248 3800 230300 3806
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223500 354 223528 3726
rect 225156 480 225184 3742
rect 225660 3726 225920 3754
rect 226764 3726 227576 3754
rect 227960 3726 228312 3754
rect 229156 3726 229416 3754
rect 230248 3742 230300 3748
rect 231032 3800 231084 3806
rect 231032 3742 231084 3748
rect 231444 3800 231496 3806
rect 231444 3742 231496 3748
rect 232228 3800 232280 3806
rect 232228 3742 232280 3748
rect 232548 3800 232600 3806
rect 232548 3742 232600 3748
rect 233424 3800 233476 3806
rect 233424 3742 233476 3748
rect 233744 3800 233796 3806
rect 233744 3742 233796 3748
rect 234620 3800 234672 3806
rect 234620 3742 234672 3748
rect 234952 3754 234980 4012
rect 236056 3754 236084 4012
rect 237252 3806 237280 4012
rect 238356 3806 238384 4012
rect 239552 3806 239580 4012
rect 240748 3806 240776 4012
rect 241852 3806 241880 4012
rect 237240 3800 237292 3806
rect 223918 354 224030 480
rect 223500 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 225892 354 225920 3726
rect 227548 480 227576 3726
rect 226310 354 226422 480
rect 225892 326 226422 354
rect 226310 -960 226422 326
rect 227506 -960 227618 480
rect 228284 354 228312 3726
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 3726
rect 231044 480 231072 3742
rect 232240 480 232268 3742
rect 233436 480 233464 3742
rect 234632 480 234660 3742
rect 234952 3726 235856 3754
rect 236056 3726 236592 3754
rect 237240 3742 237292 3748
rect 238116 3800 238168 3806
rect 238116 3742 238168 3748
rect 238344 3800 238396 3806
rect 238344 3742 238396 3748
rect 239312 3800 239364 3806
rect 239312 3742 239364 3748
rect 239540 3800 239592 3806
rect 239540 3742 239592 3748
rect 240508 3800 240560 3806
rect 240508 3742 240560 3748
rect 240736 3800 240788 3806
rect 240736 3742 240788 3748
rect 241704 3800 241756 3806
rect 241704 3742 241756 3748
rect 241840 3800 241892 3806
rect 241840 3742 241892 3748
rect 242900 3800 242952 3806
rect 242900 3742 242952 3748
rect 243048 3754 243076 4012
rect 244152 3874 244180 4012
rect 244140 3868 244192 3874
rect 244140 3810 244192 3816
rect 245200 3868 245252 3874
rect 245200 3810 245252 3816
rect 235828 480 235856 3726
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 3726
rect 238128 480 238156 3742
rect 239324 480 239352 3742
rect 240520 480 240548 3742
rect 241716 480 241744 3742
rect 242912 480 242940 3742
rect 243048 3726 244136 3754
rect 244108 480 244136 3726
rect 245212 480 245240 3810
rect 245348 3806 245376 4012
rect 246544 3806 246572 4012
rect 247648 3942 247676 4012
rect 247636 3936 247688 3942
rect 247636 3878 247688 3884
rect 248604 3936 248656 3942
rect 248604 3878 248656 3884
rect 248844 3890 248872 4012
rect 245336 3800 245388 3806
rect 245336 3742 245388 3748
rect 246396 3800 246448 3806
rect 246396 3742 246448 3748
rect 246532 3800 246584 3806
rect 246532 3742 246584 3748
rect 247592 3800 247644 3806
rect 247592 3742 247644 3748
rect 246408 480 246436 3742
rect 247604 480 247632 3742
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 236982 -960 237094 326
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248616 354 248644 3878
rect 248844 3862 248920 3890
rect 248892 2854 248920 3862
rect 250040 3806 250068 4012
rect 251144 3890 251172 4012
rect 251100 3862 251172 3890
rect 250028 3800 250080 3806
rect 250028 3742 250080 3748
rect 251100 2854 251128 3862
rect 252340 3806 252368 4012
rect 253444 3890 253472 4012
rect 254640 3890 254668 4012
rect 253400 3862 253472 3890
rect 254596 3862 254668 3890
rect 251180 3800 251232 3806
rect 251180 3742 251232 3748
rect 252328 3800 252380 3806
rect 252328 3742 252380 3748
rect 248880 2848 248932 2854
rect 248880 2790 248932 2796
rect 249984 2848 250036 2854
rect 249984 2790 250036 2796
rect 251088 2848 251140 2854
rect 251088 2790 251140 2796
rect 249996 480 250024 2790
rect 251192 480 251220 3742
rect 253400 2922 253428 3862
rect 253480 3800 253532 3806
rect 253480 3742 253532 3748
rect 253388 2916 253440 2922
rect 253388 2858 253440 2864
rect 252376 2848 252428 2854
rect 252376 2790 252428 2796
rect 252388 480 252416 2790
rect 253492 480 253520 3742
rect 254596 2854 254624 3862
rect 255836 3806 255864 4012
rect 256940 3874 256968 4012
rect 256928 3868 256980 3874
rect 256928 3810 256980 3816
rect 258136 3806 258164 4012
rect 259240 3874 259268 4012
rect 258264 3868 258316 3874
rect 258264 3810 258316 3816
rect 259228 3868 259280 3874
rect 259228 3810 259280 3816
rect 255824 3800 255876 3806
rect 255824 3742 255876 3748
rect 257068 3800 257120 3806
rect 257068 3742 257120 3748
rect 258124 3800 258176 3806
rect 258124 3742 258176 3748
rect 254676 2916 254728 2922
rect 254676 2858 254728 2864
rect 254584 2848 254636 2854
rect 254584 2790 254636 2796
rect 254688 480 254716 2858
rect 255872 2848 255924 2854
rect 255872 2790 255924 2796
rect 255884 480 255912 2790
rect 257080 480 257108 3742
rect 258276 480 258304 3810
rect 260436 3806 260464 4012
rect 261632 3874 261660 4012
rect 260656 3868 260708 3874
rect 260656 3810 260708 3816
rect 261620 3868 261672 3874
rect 261620 3810 261672 3816
rect 259460 3800 259512 3806
rect 259460 3742 259512 3748
rect 260424 3800 260476 3806
rect 260424 3742 260476 3748
rect 259472 480 259500 3742
rect 260668 480 260696 3810
rect 262736 3806 262764 4012
rect 263932 3874 263960 4012
rect 262956 3868 263008 3874
rect 262956 3810 263008 3816
rect 263920 3868 263972 3874
rect 263920 3810 263972 3816
rect 261760 3800 261812 3806
rect 261760 3742 261812 3748
rect 262724 3800 262776 3806
rect 262724 3742 262776 3748
rect 261772 480 261800 3742
rect 262968 480 262996 3810
rect 265036 3806 265064 4012
rect 265348 3868 265400 3874
rect 265348 3810 265400 3816
rect 264152 3800 264204 3806
rect 264152 3742 264204 3748
rect 265024 3800 265076 3806
rect 265024 3742 265076 3748
rect 264164 480 264192 3742
rect 265360 480 265388 3810
rect 266232 3754 266260 4012
rect 267428 3806 267456 4012
rect 268532 3874 268560 4012
rect 268520 3868 268572 3874
rect 268520 3810 268572 3816
rect 269728 3806 269756 4012
rect 270832 3874 270860 4012
rect 270040 3868 270092 3874
rect 270040 3810 270092 3816
rect 270820 3868 270872 3874
rect 270820 3810 270872 3816
rect 266544 3800 266596 3806
rect 266232 3726 266308 3754
rect 266544 3742 266596 3748
rect 267416 3800 267468 3806
rect 267416 3742 267468 3748
rect 268844 3800 268896 3806
rect 268844 3742 268896 3748
rect 269716 3800 269768 3806
rect 269716 3742 269768 3748
rect 266280 1358 266308 3726
rect 266268 1352 266320 1358
rect 266268 1294 266320 1300
rect 266556 480 266584 3742
rect 267740 1352 267792 1358
rect 267740 1294 267792 1300
rect 267752 480 267780 1294
rect 268856 480 268884 3742
rect 270052 480 270080 3810
rect 272028 3806 272056 4012
rect 272432 3868 272484 3874
rect 272432 3810 272484 3816
rect 271236 3800 271288 3806
rect 271236 3742 271288 3748
rect 272016 3800 272068 3806
rect 272016 3742 272068 3748
rect 271248 480 271276 3742
rect 272444 480 272472 3810
rect 273224 3754 273252 4012
rect 273180 3726 273252 3754
rect 273628 3800 273680 3806
rect 273628 3742 273680 3748
rect 274328 3754 274356 4012
rect 275524 3874 275552 4012
rect 275512 3868 275564 3874
rect 275512 3810 275564 3816
rect 276720 3806 276748 4012
rect 277824 3874 277852 4012
rect 277124 3868 277176 3874
rect 277124 3810 277176 3816
rect 277812 3868 277864 3874
rect 277812 3810 277864 3816
rect 276708 3800 276760 3806
rect 273180 1358 273208 3726
rect 273168 1352 273220 1358
rect 273168 1294 273220 1300
rect 273640 480 273668 3742
rect 274328 3726 274404 3754
rect 276708 3742 276760 3748
rect 274376 746 274404 3726
rect 274824 1352 274876 1358
rect 274824 1294 274876 1300
rect 274364 740 274416 746
rect 274364 682 274416 688
rect 274836 480 274864 1294
rect 276020 740 276072 746
rect 276020 682 276072 688
rect 276032 480 276060 682
rect 277136 480 277164 3810
rect 279020 3806 279048 4012
rect 279516 3868 279568 3874
rect 279516 3810 279568 3816
rect 278320 3800 278372 3806
rect 278320 3742 278372 3748
rect 279008 3800 279060 3806
rect 279008 3742 279060 3748
rect 278332 480 278360 3742
rect 279528 480 279556 3810
rect 280124 3754 280152 4012
rect 280080 3726 280152 3754
rect 280712 3800 280764 3806
rect 280712 3742 280764 3748
rect 281320 3754 281348 4012
rect 282516 3754 282544 4012
rect 283620 3806 283648 4012
rect 284816 3874 284844 4012
rect 285920 3942 285948 4012
rect 285908 3936 285960 3942
rect 285908 3878 285960 3884
rect 284804 3868 284856 3874
rect 284804 3810 284856 3816
rect 286600 3868 286652 3874
rect 286600 3810 286652 3816
rect 283608 3800 283660 3806
rect 280080 1358 280108 3726
rect 280068 1352 280120 1358
rect 280068 1294 280120 1300
rect 280724 480 280752 3742
rect 281320 3726 281396 3754
rect 282516 3726 282592 3754
rect 283608 3742 283660 3748
rect 285404 3800 285456 3806
rect 285404 3742 285456 3748
rect 281368 1290 281396 3726
rect 282564 1358 282592 3726
rect 281908 1352 281960 1358
rect 281908 1294 281960 1300
rect 282552 1352 282604 1358
rect 282552 1294 282604 1300
rect 284300 1352 284352 1358
rect 284300 1294 284352 1300
rect 281356 1284 281408 1290
rect 281356 1226 281408 1232
rect 281920 480 281948 1294
rect 283104 1284 283156 1290
rect 283104 1226 283156 1232
rect 283116 480 283144 1226
rect 284312 480 284340 1294
rect 285416 480 285444 3742
rect 286612 480 286640 3810
rect 287116 3806 287144 4012
rect 287796 3936 287848 3942
rect 287796 3878 287848 3884
rect 287104 3800 287156 3806
rect 287104 3742 287156 3748
rect 287808 480 287836 3878
rect 288312 3754 288340 4012
rect 288992 3800 289044 3806
rect 288312 3726 288388 3754
rect 288992 3742 289044 3748
rect 289416 3754 289444 4012
rect 290612 3754 290640 4012
rect 291716 3806 291744 4012
rect 292912 3874 292940 4012
rect 292900 3868 292952 3874
rect 292900 3810 292952 3816
rect 294108 3806 294136 4012
rect 294880 3868 294932 3874
rect 294880 3810 294932 3816
rect 291704 3800 291756 3806
rect 288360 1358 288388 3726
rect 288348 1352 288400 1358
rect 288348 1294 288400 1300
rect 289004 480 289032 3742
rect 289416 3726 289492 3754
rect 290612 3726 290688 3754
rect 291704 3742 291756 3748
rect 293684 3800 293736 3806
rect 293684 3742 293736 3748
rect 294096 3800 294148 3806
rect 294096 3742 294148 3748
rect 289464 1290 289492 3726
rect 290188 1352 290240 1358
rect 290188 1294 290240 1300
rect 289452 1284 289504 1290
rect 289452 1226 289504 1232
rect 290200 480 290228 1294
rect 290660 610 290688 3726
rect 291384 1284 291436 1290
rect 291384 1226 291436 1232
rect 290648 604 290700 610
rect 290648 546 290700 552
rect 291396 480 291424 1226
rect 292580 604 292632 610
rect 292580 546 292632 552
rect 292592 480 292620 546
rect 293696 480 293724 3742
rect 294892 480 294920 3810
rect 295212 3754 295240 4012
rect 296076 3800 296128 3806
rect 295212 3726 295288 3754
rect 296076 3742 296128 3748
rect 296408 3754 296436 4012
rect 297512 3754 297540 4012
rect 298708 3806 298736 4012
rect 299904 3874 299932 4012
rect 299892 3868 299944 3874
rect 299892 3810 299944 3816
rect 301008 3806 301036 4012
rect 301964 3868 302016 3874
rect 301964 3810 302016 3816
rect 298696 3800 298748 3806
rect 295260 1358 295288 3726
rect 295248 1352 295300 1358
rect 295248 1294 295300 1300
rect 296088 480 296116 3742
rect 296408 3726 296484 3754
rect 297512 3726 297588 3754
rect 298696 3742 298748 3748
rect 300768 3800 300820 3806
rect 300768 3742 300820 3748
rect 300996 3800 301048 3806
rect 300996 3742 301048 3748
rect 296456 1290 296484 3726
rect 297560 1358 297588 3726
rect 297272 1352 297324 1358
rect 297272 1294 297324 1300
rect 297548 1352 297600 1358
rect 297548 1294 297600 1300
rect 299664 1352 299716 1358
rect 299664 1294 299716 1300
rect 296444 1284 296496 1290
rect 296444 1226 296496 1232
rect 297284 480 297312 1294
rect 298468 1284 298520 1290
rect 298468 1226 298520 1232
rect 298480 480 298508 1226
rect 299676 480 299704 1294
rect 300780 480 300808 3742
rect 301976 480 302004 3810
rect 302204 3754 302232 4012
rect 302160 3726 302232 3754
rect 303160 3800 303212 3806
rect 303160 3742 303212 3748
rect 303308 3754 303336 4012
rect 304504 3754 304532 4012
rect 305700 3754 305728 4012
rect 306804 3874 306832 4012
rect 306792 3868 306844 3874
rect 306792 3810 306844 3816
rect 308000 3806 308028 4012
rect 309048 3868 309100 3874
rect 309048 3810 309100 3816
rect 307988 3800 308040 3806
rect 302160 1358 302188 3726
rect 302148 1352 302200 1358
rect 302148 1294 302200 1300
rect 303172 480 303200 3742
rect 303308 3726 303384 3754
rect 304504 3726 304580 3754
rect 305700 3726 305776 3754
rect 307988 3742 308040 3748
rect 303356 1290 303384 3726
rect 304356 1352 304408 1358
rect 304356 1294 304408 1300
rect 303344 1284 303396 1290
rect 303344 1226 303396 1232
rect 304368 480 304396 1294
rect 304552 610 304580 3726
rect 305748 1358 305776 3726
rect 305736 1352 305788 1358
rect 305736 1294 305788 1300
rect 307944 1352 307996 1358
rect 307944 1294 307996 1300
rect 305552 1284 305604 1290
rect 305552 1226 305604 1232
rect 304540 604 304592 610
rect 304540 546 304592 552
rect 305564 480 305592 1226
rect 306748 604 306800 610
rect 306748 546 306800 552
rect 306760 480 306788 546
rect 307956 480 307984 1294
rect 309060 480 309088 3810
rect 309196 3754 309224 4012
rect 310300 3890 310328 4012
rect 311496 3890 311524 4012
rect 310300 3862 310376 3890
rect 311496 3862 311572 3890
rect 310244 3800 310296 3806
rect 309196 3726 309272 3754
rect 310244 3742 310296 3748
rect 309244 2854 309272 3726
rect 309232 2848 309284 2854
rect 309232 2790 309284 2796
rect 310256 480 310284 3742
rect 310348 1358 310376 3862
rect 311440 2848 311492 2854
rect 311440 2790 311492 2796
rect 310336 1352 310388 1358
rect 310336 1294 310388 1300
rect 311452 480 311480 2790
rect 311544 1222 311572 3862
rect 312600 3754 312628 4012
rect 312556 3726 312628 3754
rect 313796 3754 313824 4012
rect 314992 3754 315020 4012
rect 316096 3806 316124 4012
rect 316084 3800 316136 3806
rect 313796 3726 313872 3754
rect 314992 3726 315068 3754
rect 317292 3754 317320 4012
rect 316084 3742 316136 3748
rect 312556 1290 312584 3726
rect 313844 1358 313872 3726
rect 315040 2854 315068 3726
rect 317248 3726 317320 3754
rect 318396 3754 318424 4012
rect 318524 3800 318576 3806
rect 318396 3726 318472 3754
rect 318524 3742 318576 3748
rect 319592 3754 319620 4012
rect 320788 3754 320816 4012
rect 321892 3754 321920 4012
rect 323088 3806 323116 4012
rect 323076 3800 323128 3806
rect 315028 2848 315080 2854
rect 315028 2790 315080 2796
rect 317248 1358 317276 3726
rect 317328 2848 317380 2854
rect 317328 2790 317380 2796
rect 312636 1352 312688 1358
rect 312636 1294 312688 1300
rect 313832 1352 313884 1358
rect 313832 1294 313884 1300
rect 316224 1352 316276 1358
rect 316224 1294 316276 1300
rect 317236 1352 317288 1358
rect 317236 1294 317288 1300
rect 312544 1284 312596 1290
rect 312544 1226 312596 1232
rect 311532 1216 311584 1222
rect 311532 1158 311584 1164
rect 312648 480 312676 1294
rect 315028 1284 315080 1290
rect 315028 1226 315080 1232
rect 313832 1216 313884 1222
rect 313832 1158 313884 1164
rect 313844 480 313872 1158
rect 315040 480 315068 1226
rect 316236 480 316264 1294
rect 317340 480 317368 2790
rect 318444 1290 318472 3726
rect 318432 1284 318484 1290
rect 318432 1226 318484 1232
rect 318536 480 318564 3742
rect 319592 3726 319668 3754
rect 320788 3726 320864 3754
rect 321892 3726 321968 3754
rect 323076 3742 323128 3748
rect 324192 3754 324220 4012
rect 325388 3754 325416 4012
rect 325608 3800 325660 3806
rect 324192 3726 324268 3754
rect 325388 3726 325464 3754
rect 325608 3742 325660 3748
rect 326584 3754 326612 4012
rect 327688 3754 327716 4012
rect 328884 3754 328912 4012
rect 329988 3754 330016 4012
rect 331184 3754 331212 4012
rect 319640 1222 319668 3726
rect 319720 1352 319772 1358
rect 319720 1294 319772 1300
rect 319628 1216 319680 1222
rect 319628 1158 319680 1164
rect 319732 480 319760 1294
rect 320836 1154 320864 3726
rect 321940 1358 321968 3726
rect 321928 1352 321980 1358
rect 321928 1294 321980 1300
rect 320916 1284 320968 1290
rect 320916 1226 320968 1232
rect 320824 1148 320876 1154
rect 320824 1090 320876 1096
rect 320928 480 320956 1226
rect 322112 1216 322164 1222
rect 322112 1158 322164 1164
rect 322124 480 322152 1158
rect 323308 1148 323360 1154
rect 323308 1090 323360 1096
rect 323320 480 323348 1090
rect 324240 610 324268 3726
rect 324412 1352 324464 1358
rect 324412 1294 324464 1300
rect 324228 604 324280 610
rect 324228 546 324280 552
rect 324424 480 324452 1294
rect 325436 1018 325464 3726
rect 325424 1012 325476 1018
rect 325424 954 325476 960
rect 325620 480 325648 3742
rect 326584 3726 326660 3754
rect 327688 3726 327764 3754
rect 328884 3726 328960 3754
rect 329988 3726 330064 3754
rect 326632 1358 326660 3726
rect 326620 1352 326672 1358
rect 326620 1294 326672 1300
rect 327736 610 327764 3726
rect 328932 1290 328960 3726
rect 329196 1352 329248 1358
rect 329196 1294 329248 1300
rect 328920 1284 328972 1290
rect 328920 1226 328972 1232
rect 328000 1012 328052 1018
rect 328000 954 328052 960
rect 326804 604 326856 610
rect 326804 546 326856 552
rect 327724 604 327776 610
rect 327724 546 327776 552
rect 326816 480 326844 546
rect 328012 480 328040 954
rect 329208 480 329236 1294
rect 330036 1222 330064 3726
rect 331140 3726 331212 3754
rect 332380 3754 332408 4012
rect 333484 3754 333512 4012
rect 334680 3754 334708 4012
rect 335876 3754 335904 4012
rect 336980 3754 337008 4012
rect 338176 3754 338204 4012
rect 339280 3754 339308 4012
rect 340476 3754 340504 4012
rect 341672 3754 341700 4012
rect 342776 3754 342804 4012
rect 343972 3754 344000 4012
rect 345076 3754 345104 4012
rect 346272 3754 346300 4012
rect 347468 3754 347496 4012
rect 348572 3754 348600 4012
rect 349768 3754 349796 4012
rect 350872 3754 350900 4012
rect 352068 3754 352096 4012
rect 353264 3754 353292 4012
rect 332380 3726 332456 3754
rect 333484 3726 333560 3754
rect 334680 3726 334756 3754
rect 335876 3726 335952 3754
rect 336980 3726 337056 3754
rect 338176 3726 338252 3754
rect 339280 3726 339356 3754
rect 340476 3726 340552 3754
rect 341672 3726 341748 3754
rect 342776 3726 342852 3754
rect 343972 3726 344048 3754
rect 345076 3726 345152 3754
rect 346272 3726 346348 3754
rect 347468 3726 347544 3754
rect 348572 3726 348648 3754
rect 349768 3726 349844 3754
rect 350872 3726 350948 3754
rect 352068 3726 352144 3754
rect 330024 1216 330076 1222
rect 330024 1158 330076 1164
rect 331140 1154 331168 3726
rect 332428 1358 332456 3726
rect 332416 1352 332468 1358
rect 332416 1294 332468 1300
rect 331588 1284 331640 1290
rect 331588 1226 331640 1232
rect 331128 1148 331180 1154
rect 331128 1090 331180 1096
rect 330392 604 330444 610
rect 330392 546 330444 552
rect 330404 480 330432 546
rect 331600 480 331628 1226
rect 332692 1216 332744 1222
rect 332692 1158 332744 1164
rect 332704 480 332732 1158
rect 333532 746 333560 3726
rect 334728 1290 334756 3726
rect 335924 1358 335952 3726
rect 335084 1352 335136 1358
rect 335084 1294 335136 1300
rect 335912 1352 335964 1358
rect 335912 1294 335964 1300
rect 334716 1284 334768 1290
rect 334716 1226 334768 1232
rect 333888 1148 333940 1154
rect 333888 1090 333940 1096
rect 333520 740 333572 746
rect 333520 682 333572 688
rect 333900 480 333928 1090
rect 335096 480 335124 1294
rect 337028 1222 337056 3726
rect 337476 1284 337528 1290
rect 337476 1226 337528 1232
rect 337016 1216 337068 1222
rect 337016 1158 337068 1164
rect 336280 740 336332 746
rect 336280 682 336332 688
rect 336292 480 336320 682
rect 337488 480 337516 1226
rect 338224 746 338252 3726
rect 339328 1358 339356 3726
rect 338672 1352 338724 1358
rect 338672 1294 338724 1300
rect 339316 1352 339368 1358
rect 339316 1294 339368 1300
rect 338212 740 338264 746
rect 338212 682 338264 688
rect 338684 480 338712 1294
rect 340524 1290 340552 3726
rect 340512 1284 340564 1290
rect 340512 1226 340564 1232
rect 341720 1222 341748 3726
rect 342168 1352 342220 1358
rect 342168 1294 342220 1300
rect 339868 1216 339920 1222
rect 339868 1158 339920 1164
rect 341708 1216 341760 1222
rect 341708 1158 341760 1164
rect 339880 480 339908 1158
rect 340972 740 341024 746
rect 340972 682 341024 688
rect 340984 480 341012 682
rect 342180 480 342208 1294
rect 342824 746 342852 3726
rect 344020 1290 344048 3726
rect 345124 1358 345152 3726
rect 345112 1352 345164 1358
rect 345112 1294 345164 1300
rect 343364 1284 343416 1290
rect 343364 1226 343416 1232
rect 344008 1284 344060 1290
rect 344008 1226 344060 1232
rect 342812 740 342864 746
rect 342812 682 342864 688
rect 343376 480 343404 1226
rect 344560 1216 344612 1222
rect 344560 1158 344612 1164
rect 344572 480 344600 1158
rect 346320 746 346348 3726
rect 346952 1284 347004 1290
rect 346952 1226 347004 1232
rect 345756 740 345808 746
rect 345756 682 345808 688
rect 346308 740 346360 746
rect 346308 682 346360 688
rect 345768 480 345796 682
rect 346964 480 346992 1226
rect 347516 882 347544 3726
rect 348056 1352 348108 1358
rect 348056 1294 348108 1300
rect 347504 876 347556 882
rect 347504 818 347556 824
rect 348068 480 348096 1294
rect 348620 1290 348648 3726
rect 349816 1358 349844 3726
rect 349804 1352 349856 1358
rect 349804 1294 349856 1300
rect 348608 1284 348660 1290
rect 348608 1226 348660 1232
rect 350448 876 350500 882
rect 350448 818 350500 824
rect 349252 740 349304 746
rect 349252 682 349304 688
rect 349264 480 349292 682
rect 350460 480 350488 818
rect 350920 746 350948 3726
rect 352116 1290 352144 3726
rect 353220 3726 353292 3754
rect 354368 3754 354396 4012
rect 355564 3754 355592 4012
rect 356668 3754 356696 4012
rect 357864 3754 357892 4012
rect 359060 3754 359088 4012
rect 360164 3754 360192 4012
rect 354368 3726 354444 3754
rect 355564 3726 355640 3754
rect 356668 3726 356744 3754
rect 357864 3726 357940 3754
rect 359060 3726 359136 3754
rect 353220 1358 353248 3726
rect 352840 1352 352892 1358
rect 352840 1294 352892 1300
rect 353208 1352 353260 1358
rect 353208 1294 353260 1300
rect 351644 1284 351696 1290
rect 351644 1226 351696 1232
rect 352104 1284 352156 1290
rect 352104 1226 352156 1232
rect 350908 740 350960 746
rect 350908 682 350960 688
rect 351656 480 351684 1226
rect 352852 480 352880 1294
rect 354036 740 354088 746
rect 354036 682 354088 688
rect 354048 480 354076 682
rect 248758 354 248870 480
rect 248616 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 354416 66 354444 3726
rect 355612 1290 355640 3726
rect 356716 1358 356744 3726
rect 356336 1352 356388 1358
rect 356336 1294 356388 1300
rect 356704 1352 356756 1358
rect 356704 1294 356756 1300
rect 355232 1284 355284 1290
rect 355232 1226 355284 1232
rect 355600 1284 355652 1290
rect 355600 1226 355652 1232
rect 355244 480 355272 1226
rect 356348 480 356376 1294
rect 357912 1222 357940 3726
rect 359108 1290 359136 3726
rect 360120 3726 360192 3754
rect 361360 3754 361388 4012
rect 362556 3754 362584 4012
rect 363660 3754 363688 4012
rect 364856 3754 364884 4012
rect 365960 3754 365988 4012
rect 367156 3754 367184 4012
rect 368352 3754 368380 4012
rect 369456 3754 369484 4012
rect 370652 3754 370680 4012
rect 371756 3754 371784 4012
rect 372952 3754 372980 4012
rect 374148 3754 374176 4012
rect 375252 3754 375280 4012
rect 376448 3754 376476 4012
rect 361360 3726 361436 3754
rect 362556 3726 362632 3754
rect 363660 3726 363736 3754
rect 364856 3726 364932 3754
rect 365960 3726 366036 3754
rect 367156 3726 367232 3754
rect 368352 3726 368428 3754
rect 369456 3726 369532 3754
rect 370652 3726 370728 3754
rect 371756 3726 371832 3754
rect 372952 3726 373028 3754
rect 374148 3726 374224 3754
rect 375252 3726 375328 3754
rect 359924 1352 359976 1358
rect 359924 1294 359976 1300
rect 358728 1284 358780 1290
rect 358728 1226 358780 1232
rect 359096 1284 359148 1290
rect 359096 1226 359148 1232
rect 357900 1216 357952 1222
rect 357900 1158 357952 1164
rect 358740 480 358768 1226
rect 359936 480 359964 1294
rect 360120 1154 360148 3726
rect 361120 1216 361172 1222
rect 361120 1158 361172 1164
rect 360108 1148 360160 1154
rect 360108 1090 360160 1096
rect 361132 480 361160 1158
rect 361408 882 361436 3726
rect 362604 1358 362632 3726
rect 362592 1352 362644 1358
rect 362592 1294 362644 1300
rect 363708 1290 363736 3726
rect 362316 1284 362368 1290
rect 362316 1226 362368 1232
rect 363696 1284 363748 1290
rect 363696 1226 363748 1232
rect 361396 876 361448 882
rect 361396 818 361448 824
rect 362328 480 362356 1226
rect 364904 1222 364932 3726
rect 365812 1352 365864 1358
rect 365812 1294 365864 1300
rect 364892 1216 364944 1222
rect 364892 1158 364944 1164
rect 363512 1148 363564 1154
rect 363512 1090 363564 1096
rect 363524 480 363552 1090
rect 364616 876 364668 882
rect 364616 818 364668 824
rect 364628 480 364656 818
rect 365824 480 365852 1294
rect 366008 746 366036 3726
rect 367204 1358 367232 3726
rect 367192 1352 367244 1358
rect 367192 1294 367244 1300
rect 367008 1284 367060 1290
rect 367008 1226 367060 1232
rect 365996 740 366048 746
rect 365996 682 366048 688
rect 367020 480 367048 1226
rect 368204 1216 368256 1222
rect 368204 1158 368256 1164
rect 368216 480 368244 1158
rect 368400 882 368428 3726
rect 368388 876 368440 882
rect 368388 818 368440 824
rect 369504 746 369532 3726
rect 370700 1358 370728 3726
rect 370596 1352 370648 1358
rect 370596 1294 370648 1300
rect 370688 1352 370740 1358
rect 370688 1294 370740 1300
rect 369400 740 369452 746
rect 369400 682 369452 688
rect 369492 740 369544 746
rect 369492 682 369544 688
rect 369412 480 369440 682
rect 370608 480 370636 1294
rect 371804 882 371832 3726
rect 373000 1290 373028 3726
rect 374092 1352 374144 1358
rect 374092 1294 374144 1300
rect 372988 1284 373040 1290
rect 372988 1226 373040 1232
rect 371700 876 371752 882
rect 371700 818 371752 824
rect 371792 876 371844 882
rect 371792 818 371844 824
rect 371712 480 371740 818
rect 372896 740 372948 746
rect 372896 682 372948 688
rect 372908 480 372936 682
rect 374104 480 374132 1294
rect 374196 1018 374224 3726
rect 375300 1222 375328 3726
rect 376404 3726 376476 3754
rect 377552 3754 377580 4012
rect 378748 3754 378776 4012
rect 379944 3754 379972 4012
rect 377552 3726 377628 3754
rect 378748 3726 378824 3754
rect 376404 1358 376432 3726
rect 376392 1352 376444 1358
rect 376392 1294 376444 1300
rect 377600 1290 377628 3726
rect 376484 1284 376536 1290
rect 376484 1226 376536 1232
rect 377588 1284 377640 1290
rect 377588 1226 377640 1232
rect 375288 1216 375340 1222
rect 375288 1158 375340 1164
rect 374184 1012 374236 1018
rect 374184 954 374236 960
rect 375288 876 375340 882
rect 375288 818 375340 824
rect 375300 480 375328 818
rect 376496 480 376524 1226
rect 378796 1086 378824 3726
rect 379900 3726 379972 3754
rect 381048 3754 381076 4012
rect 382244 3754 382272 4012
rect 381048 3726 381124 3754
rect 378876 1216 378928 1222
rect 378876 1158 378928 1164
rect 378784 1080 378836 1086
rect 378784 1022 378836 1028
rect 377680 1012 377732 1018
rect 377680 954 377732 960
rect 377692 480 377720 954
rect 378888 480 378916 1158
rect 379900 1018 379928 3726
rect 379980 1352 380032 1358
rect 379980 1294 380032 1300
rect 379888 1012 379940 1018
rect 379888 954 379940 960
rect 379992 480 380020 1294
rect 381096 1222 381124 3726
rect 382200 3726 382272 3754
rect 383348 3754 383376 4012
rect 384544 3754 384572 4012
rect 385740 3754 385768 4012
rect 386844 3754 386872 4012
rect 388040 3754 388068 4012
rect 389236 3754 389264 4012
rect 390340 3754 390368 4012
rect 391536 3754 391564 4012
rect 392640 3754 392668 4012
rect 393836 3754 393864 4012
rect 395032 3754 395060 4012
rect 396136 3754 396164 4012
rect 397332 3754 397360 4012
rect 398436 3754 398464 4012
rect 399632 3754 399660 4012
rect 400828 3754 400856 4012
rect 401932 3754 401960 4012
rect 403128 3754 403156 4012
rect 404232 3754 404260 4012
rect 405428 3754 405456 4012
rect 406624 3754 406652 4012
rect 407728 3754 407756 4012
rect 408924 3754 408952 4012
rect 410028 3754 410056 4012
rect 411224 3754 411252 4012
rect 383348 3726 383424 3754
rect 384544 3726 384620 3754
rect 385740 3726 385816 3754
rect 386844 3726 386920 3754
rect 388040 3726 388116 3754
rect 389236 3726 389312 3754
rect 390340 3726 390416 3754
rect 391536 3726 391612 3754
rect 392640 3726 392716 3754
rect 393836 3726 393912 3754
rect 395032 3726 395108 3754
rect 396136 3726 396212 3754
rect 397332 3726 397408 3754
rect 398436 3726 398512 3754
rect 399632 3726 399708 3754
rect 400828 3726 400904 3754
rect 401932 3726 402008 3754
rect 403128 3726 403204 3754
rect 404232 3726 404308 3754
rect 405428 3726 405504 3754
rect 406624 3726 406700 3754
rect 407728 3726 407804 3754
rect 408924 3726 409000 3754
rect 410028 3726 410104 3754
rect 381176 1284 381228 1290
rect 381176 1226 381228 1232
rect 381084 1216 381136 1222
rect 381084 1158 381136 1164
rect 381188 480 381216 1226
rect 382200 1154 382228 3726
rect 382188 1148 382240 1154
rect 382188 1090 382240 1096
rect 382372 1080 382424 1086
rect 382372 1022 382424 1028
rect 382384 480 382412 1022
rect 354404 60 354456 66
rect 354404 2 354456 8
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 82 357614 480
rect 357360 66 357614 82
rect 357348 60 357614 66
rect 357400 54 357614 60
rect 357348 2 357400 8
rect 357502 -960 357614 54
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383396 338 383424 3726
rect 383568 1012 383620 1018
rect 383568 954 383620 960
rect 383580 480 383608 954
rect 384592 882 384620 3726
rect 385788 1358 385816 3726
rect 385776 1352 385828 1358
rect 385776 1294 385828 1300
rect 384764 1216 384816 1222
rect 384764 1158 384816 1164
rect 384580 876 384632 882
rect 384580 818 384632 824
rect 384776 480 384804 1158
rect 385960 1148 386012 1154
rect 385960 1090 386012 1096
rect 385972 480 386000 1090
rect 386892 1086 386920 3726
rect 388088 1290 388116 3726
rect 388076 1284 388128 1290
rect 388076 1226 388128 1232
rect 389284 1154 389312 3726
rect 389456 1352 389508 1358
rect 389456 1294 389508 1300
rect 389272 1148 389324 1154
rect 389272 1090 389324 1096
rect 386880 1080 386932 1086
rect 386880 1022 386932 1028
rect 388260 876 388312 882
rect 388260 818 388312 824
rect 388272 480 388300 818
rect 389468 480 389496 1294
rect 390388 1222 390416 3726
rect 390376 1216 390428 1222
rect 390376 1158 390428 1164
rect 390652 1080 390704 1086
rect 390652 1022 390704 1028
rect 390664 480 390692 1022
rect 391584 882 391612 3726
rect 391848 1284 391900 1290
rect 391848 1226 391900 1232
rect 391572 876 391624 882
rect 391572 818 391624 824
rect 391860 480 391888 1226
rect 383384 332 383436 338
rect 383384 274 383436 280
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 354 387238 480
rect 386800 338 387238 354
rect 386788 332 387238 338
rect 386840 326 387238 332
rect 386788 274 386840 280
rect 387126 -960 387238 326
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392688 134 392716 3726
rect 393884 1290 393912 3726
rect 395080 1358 395108 3726
rect 395068 1352 395120 1358
rect 395068 1294 395120 1300
rect 393872 1284 393924 1290
rect 393872 1226 393924 1232
rect 396184 1222 396212 3726
rect 394240 1216 394292 1222
rect 394240 1158 394292 1164
rect 396172 1216 396224 1222
rect 396172 1158 396224 1164
rect 393044 1148 393096 1154
rect 393044 1090 393096 1096
rect 393056 480 393084 1090
rect 394252 480 394280 1158
rect 397380 882 397408 3726
rect 397736 1284 397788 1290
rect 397736 1226 397788 1232
rect 395344 876 395396 882
rect 395344 818 395396 824
rect 397368 876 397420 882
rect 397368 818 397420 824
rect 395356 480 395384 818
rect 397748 480 397776 1226
rect 398484 1154 398512 3726
rect 399680 1358 399708 3726
rect 398932 1352 398984 1358
rect 398932 1294 398984 1300
rect 399668 1352 399720 1358
rect 399668 1294 399720 1300
rect 398472 1148 398524 1154
rect 398472 1090 398524 1096
rect 398944 480 398972 1294
rect 400876 1222 400904 3726
rect 400128 1216 400180 1222
rect 400128 1158 400180 1164
rect 400864 1216 400916 1222
rect 400864 1158 400916 1164
rect 400140 480 400168 1158
rect 401324 876 401376 882
rect 401324 818 401376 824
rect 401336 480 401364 818
rect 392676 128 392728 134
rect 392676 70 392728 76
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396172 128 396224 134
rect 396510 82 396622 480
rect 396224 76 396622 82
rect 396172 70 396622 76
rect 396184 54 396622 70
rect 396510 -960 396622 54
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 401980 134 402008 3726
rect 403176 1290 403204 3726
rect 403624 1352 403676 1358
rect 403624 1294 403676 1300
rect 403164 1284 403216 1290
rect 403164 1226 403216 1232
rect 402520 1148 402572 1154
rect 402520 1090 402572 1096
rect 402532 480 402560 1090
rect 403636 480 403664 1294
rect 404280 1154 404308 3726
rect 405476 1358 405504 3726
rect 405464 1352 405516 1358
rect 405464 1294 405516 1300
rect 404820 1216 404872 1222
rect 404820 1158 404872 1164
rect 404268 1148 404320 1154
rect 404268 1090 404320 1096
rect 404832 480 404860 1158
rect 406672 882 406700 3726
rect 407212 1284 407264 1290
rect 407212 1226 407264 1232
rect 406660 876 406712 882
rect 406660 818 406712 824
rect 407224 480 407252 1226
rect 407776 1222 407804 3726
rect 407764 1216 407816 1222
rect 407764 1158 407816 1164
rect 408972 1154 409000 3726
rect 409604 1352 409656 1358
rect 409604 1294 409656 1300
rect 408408 1148 408460 1154
rect 408408 1090 408460 1096
rect 408960 1148 409012 1154
rect 408960 1090 409012 1096
rect 408420 480 408448 1090
rect 409616 480 409644 1294
rect 410076 1290 410104 3726
rect 411180 3726 411252 3754
rect 412420 3754 412448 4012
rect 413524 3754 413552 4012
rect 414720 3754 414748 4012
rect 415916 3754 415944 4012
rect 417020 3754 417048 4012
rect 418216 3754 418244 4012
rect 419320 3754 419348 4012
rect 420516 3754 420544 4012
rect 421712 3754 421740 4012
rect 422816 3754 422844 4012
rect 424012 3754 424040 4012
rect 425116 3754 425144 4012
rect 426312 3754 426340 4012
rect 427508 3754 427536 4012
rect 428612 3754 428640 4012
rect 429808 3754 429836 4012
rect 430912 3754 430940 4012
rect 432108 3754 432136 4012
rect 433304 3754 433332 4012
rect 434408 3754 434436 4012
rect 412420 3726 412496 3754
rect 413524 3726 413600 3754
rect 414720 3726 414796 3754
rect 415916 3726 415992 3754
rect 417020 3726 417096 3754
rect 418216 3726 418292 3754
rect 419320 3726 419396 3754
rect 420516 3726 420592 3754
rect 421712 3726 421788 3754
rect 422816 3726 422892 3754
rect 424012 3726 424088 3754
rect 425116 3726 425192 3754
rect 426312 3726 426388 3754
rect 427508 3726 427584 3754
rect 428612 3726 428688 3754
rect 429808 3726 429884 3754
rect 430912 3726 431080 3754
rect 432108 3726 432184 3754
rect 411180 2854 411208 3726
rect 411168 2848 411220 2854
rect 411168 2790 411220 2796
rect 410064 1284 410116 1290
rect 410064 1226 410116 1232
rect 411904 1216 411956 1222
rect 411904 1158 411956 1164
rect 410800 876 410852 882
rect 410800 818 410852 824
rect 410812 480 410840 818
rect 411916 480 411944 1158
rect 401968 128 402020 134
rect 401968 70 402020 76
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 82 406098 480
rect 406200 128 406252 134
rect 405986 76 406200 82
rect 405986 70 406252 76
rect 405986 54 406240 70
rect 405986 -960 406098 54
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412468 202 412496 3726
rect 413572 1358 413600 3726
rect 413560 1352 413612 1358
rect 413560 1294 413612 1300
rect 414296 1284 414348 1290
rect 414296 1226 414348 1232
rect 413100 1148 413152 1154
rect 413100 1090 413152 1096
rect 413112 480 413140 1090
rect 414308 480 414336 1226
rect 414768 1018 414796 3726
rect 415492 2848 415544 2854
rect 415492 2790 415544 2796
rect 414756 1012 414808 1018
rect 414756 954 414808 960
rect 415504 480 415532 2790
rect 415964 1154 415992 3726
rect 415952 1148 416004 1154
rect 415952 1090 416004 1096
rect 417068 1086 417096 3726
rect 417884 1352 417936 1358
rect 417884 1294 417936 1300
rect 417056 1080 417108 1086
rect 417056 1022 417108 1028
rect 417896 480 417924 1294
rect 418264 1290 418292 3726
rect 418252 1284 418304 1290
rect 418252 1226 418304 1232
rect 418988 1012 419040 1018
rect 418988 954 419040 960
rect 419000 480 419028 954
rect 419368 882 419396 3726
rect 420564 1222 420592 3726
rect 420552 1216 420604 1222
rect 420552 1158 420604 1164
rect 420184 1148 420236 1154
rect 420184 1090 420236 1096
rect 419356 876 419408 882
rect 419356 818 419408 824
rect 420196 480 420224 1090
rect 421380 1080 421432 1086
rect 421380 1022 421432 1028
rect 421392 480 421420 1022
rect 412456 196 412508 202
rect 412456 138 412508 144
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 218 416770 480
rect 416658 202 416912 218
rect 416658 196 416924 202
rect 416658 190 416872 196
rect 416658 -960 416770 190
rect 416872 138 416924 144
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 421760 134 421788 3726
rect 422864 1358 422892 3726
rect 422852 1352 422904 1358
rect 422852 1294 422904 1300
rect 422576 1284 422628 1290
rect 422576 1226 422628 1232
rect 422588 480 422616 1226
rect 424060 1018 424088 3726
rect 425164 1222 425192 3726
rect 426360 1290 426388 3726
rect 427556 1358 427584 3726
rect 427268 1352 427320 1358
rect 427268 1294 427320 1300
rect 427544 1352 427596 1358
rect 427544 1294 427596 1300
rect 426348 1284 426400 1290
rect 426348 1226 426400 1232
rect 424968 1216 425020 1222
rect 424968 1158 425020 1164
rect 425152 1216 425204 1222
rect 425152 1158 425204 1164
rect 424048 1012 424100 1018
rect 424048 954 424100 960
rect 423404 876 423456 882
rect 423404 818 423456 824
rect 421748 128 421800 134
rect 421748 70 421800 76
rect 422546 -960 422658 480
rect 423416 354 423444 818
rect 424980 480 425008 1158
rect 427280 480 427308 1294
rect 428660 1154 428688 3726
rect 429660 1216 429712 1222
rect 429660 1158 429712 1164
rect 428648 1148 428700 1154
rect 428648 1090 428700 1096
rect 428464 1012 428516 1018
rect 428464 954 428516 960
rect 428476 480 428504 954
rect 429672 480 429700 1158
rect 429856 882 429884 3726
rect 430856 1284 430908 1290
rect 430856 1226 430908 1232
rect 429844 876 429896 882
rect 429844 818 429896 824
rect 430868 480 430896 1226
rect 423742 354 423854 480
rect 423416 326 423854 354
rect 423742 -960 423854 326
rect 424938 -960 425050 480
rect 425796 128 425848 134
rect 426134 82 426246 480
rect 425848 76 426246 82
rect 425796 70 426246 76
rect 425808 54 426246 70
rect 426134 -960 426246 54
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 431052 134 431080 3726
rect 431868 1352 431920 1358
rect 431868 1294 431920 1300
rect 431880 354 431908 1294
rect 432156 1018 432184 3726
rect 433260 3726 433332 3754
rect 434364 3726 434436 3754
rect 435604 3754 435632 4012
rect 436708 3754 436736 4012
rect 437904 3754 437932 4012
rect 439100 3754 439128 4012
rect 440204 3754 440232 4012
rect 435604 3726 435680 3754
rect 436708 3726 436784 3754
rect 437904 3726 437980 3754
rect 439100 3726 439176 3754
rect 433260 1358 433288 3726
rect 433248 1352 433300 1358
rect 433248 1294 433300 1300
rect 433248 1148 433300 1154
rect 433248 1090 433300 1096
rect 432144 1012 432196 1018
rect 432144 954 432196 960
rect 433260 480 433288 1090
rect 434364 950 434392 3726
rect 435652 1290 435680 3726
rect 435640 1284 435692 1290
rect 435640 1226 435692 1232
rect 436756 1222 436784 3726
rect 437848 1352 437900 1358
rect 437848 1294 437900 1300
rect 436744 1216 436796 1222
rect 436744 1158 436796 1164
rect 436744 1012 436796 1018
rect 436744 954 436796 960
rect 434352 944 434404 950
rect 434352 886 434404 892
rect 434444 876 434496 882
rect 434444 818 434496 824
rect 434456 480 434484 818
rect 436756 480 436784 954
rect 437860 898 437888 1294
rect 437952 1086 437980 3726
rect 439148 1154 439176 3726
rect 440160 3726 440232 3754
rect 441400 3754 441428 4012
rect 442596 3754 442624 4012
rect 443700 3754 443728 4012
rect 444896 3754 444924 4012
rect 446000 3754 446028 4012
rect 447196 3754 447224 4012
rect 448392 3754 448420 4012
rect 449496 3754 449524 4012
rect 450692 3754 450720 4012
rect 451796 3754 451824 4012
rect 452992 3754 453020 4012
rect 454188 3754 454216 4012
rect 455292 3754 455320 4012
rect 456488 3754 456516 4012
rect 457592 3754 457620 4012
rect 458788 3754 458816 4012
rect 459984 3754 460012 4012
rect 461088 3754 461116 4012
rect 462284 3754 462312 4012
rect 441400 3726 441476 3754
rect 442596 3726 442672 3754
rect 443700 3726 443776 3754
rect 444896 3726 444972 3754
rect 446000 3726 446076 3754
rect 447196 3726 447272 3754
rect 448392 3726 448468 3754
rect 449496 3726 449572 3754
rect 450692 3726 450768 3754
rect 451796 3726 451872 3754
rect 452992 3726 453068 3754
rect 454188 3726 454264 3754
rect 455292 3726 455368 3754
rect 456488 3726 456564 3754
rect 457592 3726 457668 3754
rect 458788 3726 458864 3754
rect 459984 3726 460060 3754
rect 461088 3726 461164 3754
rect 440160 2854 440188 3726
rect 440148 2848 440200 2854
rect 440148 2790 440200 2796
rect 441448 1358 441476 3726
rect 441436 1352 441488 1358
rect 441436 1294 441488 1300
rect 442644 1290 442672 3726
rect 439964 1284 440016 1290
rect 439964 1226 440016 1232
rect 442632 1284 442684 1290
rect 442632 1226 442684 1232
rect 439136 1148 439188 1154
rect 439136 1090 439188 1096
rect 437940 1080 437992 1086
rect 437940 1022 437992 1028
rect 439136 944 439188 950
rect 437860 870 437980 898
rect 439136 886 439188 892
rect 437952 480 437980 870
rect 439148 480 439176 886
rect 432022 354 432134 480
rect 431880 326 432134 354
rect 431040 128 431092 134
rect 431040 70 431092 76
rect 432022 -960 432134 326
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435180 128 435232 134
rect 435518 82 435630 480
rect 435232 76 435630 82
rect 435180 70 435630 76
rect 435192 54 435630 70
rect 435518 -960 435630 54
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 439976 354 440004 1226
rect 441528 1216 441580 1222
rect 441528 1158 441580 1164
rect 441540 480 441568 1158
rect 442632 1080 442684 1086
rect 442632 1022 442684 1028
rect 442644 480 442672 1022
rect 443748 882 443776 3726
rect 444944 1222 444972 3726
rect 445024 2848 445076 2854
rect 445024 2790 445076 2796
rect 444932 1216 444984 1222
rect 444932 1158 444984 1164
rect 443828 1148 443880 1154
rect 443828 1090 443880 1096
rect 443736 876 443788 882
rect 443736 818 443788 824
rect 443840 480 443868 1090
rect 445036 480 445064 2790
rect 445852 1352 445904 1358
rect 445852 1294 445904 1300
rect 440302 354 440414 480
rect 439976 326 440414 354
rect 440302 -960 440414 326
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445864 354 445892 1294
rect 446048 1086 446076 3726
rect 447244 1358 447272 3726
rect 447232 1352 447284 1358
rect 447232 1294 447284 1300
rect 447416 1284 447468 1290
rect 447416 1226 447468 1232
rect 446036 1080 446088 1086
rect 446036 1022 446088 1028
rect 447428 480 447456 1226
rect 448440 1154 448468 3726
rect 449544 2854 449572 3726
rect 449532 2848 449584 2854
rect 449532 2790 449584 2796
rect 450740 1222 450768 3726
rect 449808 1216 449860 1222
rect 449808 1158 449860 1164
rect 450728 1216 450780 1222
rect 450728 1158 450780 1164
rect 448428 1148 448480 1154
rect 448428 1090 448480 1096
rect 448244 876 448296 882
rect 448244 818 448296 824
rect 446190 354 446302 480
rect 445864 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448256 354 448284 818
rect 449820 480 449848 1158
rect 450912 1080 450964 1086
rect 450912 1022 450964 1028
rect 450924 480 450952 1022
rect 451844 882 451872 3726
rect 453040 1358 453068 3726
rect 452108 1352 452160 1358
rect 452108 1294 452160 1300
rect 453028 1352 453080 1358
rect 453028 1294 453080 1300
rect 451832 876 451884 882
rect 451832 818 451884 824
rect 452120 480 452148 1294
rect 454236 1154 454264 3726
rect 454500 2848 454552 2854
rect 454500 2790 454552 2796
rect 453304 1148 453356 1154
rect 453304 1090 453356 1096
rect 454224 1148 454276 1154
rect 454224 1090 454276 1096
rect 453316 480 453344 1090
rect 454512 480 454540 2790
rect 455340 1086 455368 3726
rect 456536 1222 456564 3726
rect 457640 1290 457668 3726
rect 458836 1358 458864 3726
rect 458088 1352 458140 1358
rect 458088 1294 458140 1300
rect 458824 1352 458876 1358
rect 458824 1294 458876 1300
rect 457628 1284 457680 1290
rect 457628 1226 457680 1232
rect 455696 1216 455748 1222
rect 455696 1158 455748 1164
rect 456524 1216 456576 1222
rect 456524 1158 456576 1164
rect 455328 1080 455380 1086
rect 455328 1022 455380 1028
rect 455708 480 455736 1158
rect 456524 876 456576 882
rect 456524 818 456576 824
rect 448582 354 448694 480
rect 448256 326 448694 354
rect 448582 -960 448694 326
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456536 354 456564 818
rect 458100 480 458128 1294
rect 459192 1148 459244 1154
rect 459192 1090 459244 1096
rect 459204 480 459232 1090
rect 456862 354 456974 480
rect 456536 326 456974 354
rect 456862 -960 456974 326
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460032 134 460060 3726
rect 461136 1086 461164 3726
rect 462240 3726 462312 3754
rect 463388 3754 463416 4012
rect 464584 3754 464612 4012
rect 465780 3754 465808 4012
rect 466884 3754 466912 4012
rect 468080 3754 468108 4012
rect 469276 3754 469304 4012
rect 470380 3754 470408 4012
rect 471576 3754 471604 4012
rect 472680 3754 472708 4012
rect 473876 3754 473904 4012
rect 475072 3754 475100 4012
rect 476176 3754 476204 4012
rect 477372 3754 477400 4012
rect 478476 3754 478504 4012
rect 479672 3754 479700 4012
rect 480868 3754 480896 4012
rect 481972 3754 482000 4012
rect 483168 3754 483196 4012
rect 484272 3754 484300 4012
rect 485468 3754 485496 4012
rect 486664 3754 486692 4012
rect 487768 3754 487796 4012
rect 488964 3754 488992 4012
rect 490068 3754 490096 4012
rect 491264 3754 491292 4012
rect 463388 3726 463464 3754
rect 464584 3726 464660 3754
rect 465780 3726 465856 3754
rect 466884 3726 466960 3754
rect 468080 3726 468156 3754
rect 469276 3726 469352 3754
rect 470380 3726 470456 3754
rect 471576 3726 471652 3754
rect 472680 3726 472756 3754
rect 473876 3726 473952 3754
rect 475072 3726 475148 3754
rect 476176 3726 476252 3754
rect 477372 3726 477448 3754
rect 478476 3726 478552 3754
rect 479672 3726 479748 3754
rect 480868 3726 480944 3754
rect 481972 3726 482048 3754
rect 483168 3726 483244 3754
rect 484272 3726 484348 3754
rect 485468 3726 485544 3754
rect 486664 3726 486740 3754
rect 487768 3726 487844 3754
rect 488964 3726 489040 3754
rect 490068 3726 490144 3754
rect 462240 1222 462268 3726
rect 462412 1284 462464 1290
rect 462412 1226 462464 1232
rect 461584 1216 461636 1222
rect 461584 1158 461636 1164
rect 462228 1216 462280 1222
rect 462228 1158 462280 1164
rect 460112 1080 460164 1086
rect 460112 1022 460164 1028
rect 461124 1080 461176 1086
rect 461124 1022 461176 1028
rect 460124 354 460152 1022
rect 461596 480 461624 1158
rect 460358 354 460470 480
rect 460124 326 460470 354
rect 460020 128 460072 134
rect 460020 70 460072 76
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462424 354 462452 1226
rect 463436 950 463464 3726
rect 463976 1352 464028 1358
rect 463976 1294 464028 1300
rect 463424 944 463476 950
rect 463424 886 463476 892
rect 463988 480 464016 1294
rect 464632 1018 464660 3726
rect 465828 1154 465856 3726
rect 465816 1148 465868 1154
rect 465816 1090 465868 1096
rect 466932 1086 466960 3726
rect 468128 1290 468156 3726
rect 468116 1284 468168 1290
rect 468116 1226 468168 1232
rect 467472 1216 467524 1222
rect 467472 1158 467524 1164
rect 466276 1080 466328 1086
rect 466276 1022 466328 1028
rect 466920 1080 466972 1086
rect 466920 1022 466972 1028
rect 464620 1012 464672 1018
rect 464620 954 464672 960
rect 466288 480 466316 1022
rect 467484 480 467512 1158
rect 468668 944 468720 950
rect 468668 886 468720 892
rect 468680 480 468708 886
rect 462750 354 462862 480
rect 462424 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 464988 128 465040 134
rect 465142 82 465254 480
rect 465040 76 465254 82
rect 464988 70 465254 76
rect 465000 54 465254 70
rect 465142 -960 465254 54
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469324 270 469352 3726
rect 469864 1012 469916 1018
rect 469864 954 469916 960
rect 469876 480 469904 954
rect 469312 264 469364 270
rect 469312 206 469364 212
rect 469834 -960 469946 480
rect 470428 202 470456 3726
rect 471624 1358 471652 3726
rect 471612 1352 471664 1358
rect 471612 1294 471664 1300
rect 472728 1222 472756 3726
rect 473084 1284 473136 1290
rect 473084 1226 473136 1232
rect 472716 1216 472768 1222
rect 472716 1158 472768 1164
rect 470692 1148 470744 1154
rect 470692 1090 470744 1096
rect 470704 354 470732 1090
rect 472256 1080 472308 1086
rect 472256 1022 472308 1028
rect 472268 480 472296 1022
rect 471030 354 471142 480
rect 470704 326 471142 354
rect 470416 196 470468 202
rect 470416 138 470468 144
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473096 354 473124 1226
rect 473924 1018 473952 3726
rect 475120 1290 475148 3726
rect 475108 1284 475160 1290
rect 475108 1226 475160 1232
rect 473912 1012 473964 1018
rect 473912 954 473964 960
rect 476224 882 476252 3726
rect 477420 1358 477448 3726
rect 478524 2854 478552 3726
rect 478512 2848 478564 2854
rect 478512 2790 478564 2796
rect 476580 1352 476632 1358
rect 476580 1294 476632 1300
rect 477408 1352 477460 1358
rect 477408 1294 477460 1300
rect 476212 876 476264 882
rect 476212 818 476264 824
rect 473422 354 473534 480
rect 473096 326 473534 354
rect 473422 -960 473534 326
rect 474188 264 474240 270
rect 474526 218 474638 480
rect 474240 212 474638 218
rect 474188 206 474638 212
rect 474200 190 474638 206
rect 474526 -960 474638 190
rect 475722 218 475834 480
rect 476592 354 476620 1294
rect 478144 1216 478196 1222
rect 478144 1158 478196 1164
rect 478156 480 478184 1158
rect 479720 1086 479748 3726
rect 480536 1284 480588 1290
rect 480536 1226 480588 1232
rect 479708 1080 479760 1086
rect 479708 1022 479760 1028
rect 479340 1012 479392 1018
rect 479340 954 479392 960
rect 479352 480 479380 954
rect 480548 480 480576 1226
rect 480916 1222 480944 3726
rect 480904 1216 480956 1222
rect 480904 1158 480956 1164
rect 482020 1154 482048 3726
rect 483216 1358 483244 3726
rect 484032 2848 484084 2854
rect 484032 2790 484084 2796
rect 482468 1352 482520 1358
rect 482468 1294 482520 1300
rect 483204 1352 483256 1358
rect 483204 1294 483256 1300
rect 482008 1148 482060 1154
rect 482008 1090 482060 1096
rect 481364 876 481416 882
rect 481364 818 481416 824
rect 476918 354 477030 480
rect 476592 326 477030 354
rect 475722 202 475976 218
rect 475722 196 475988 202
rect 475722 190 475936 196
rect 475722 -960 475834 190
rect 475936 138 475988 144
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481376 354 481404 818
rect 481702 354 481814 480
rect 481376 326 481814 354
rect 482480 354 482508 1294
rect 484044 480 484072 2790
rect 484320 950 484348 3726
rect 485516 1290 485544 3726
rect 485504 1284 485556 1290
rect 485504 1226 485556 1232
rect 486712 1222 486740 3726
rect 487816 2854 487844 3726
rect 487804 2848 487856 2854
rect 487804 2790 487856 2796
rect 488816 1352 488868 1358
rect 488816 1294 488868 1300
rect 486424 1216 486476 1222
rect 486424 1158 486476 1164
rect 486700 1216 486752 1222
rect 486700 1158 486752 1164
rect 484860 1080 484912 1086
rect 484860 1022 484912 1028
rect 484308 944 484360 950
rect 484308 886 484360 892
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 481702 -960 481814 326
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484872 354 484900 1022
rect 486436 480 486464 1158
rect 487252 1148 487304 1154
rect 487252 1090 487304 1096
rect 485198 354 485310 480
rect 484872 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487264 354 487292 1090
rect 488828 480 488856 1294
rect 489012 1154 489040 3726
rect 490116 1358 490144 3726
rect 491220 3726 491292 3754
rect 492460 3754 492488 4012
rect 493564 3754 493592 4012
rect 494760 3754 494788 4012
rect 495956 3754 495984 4012
rect 497060 3754 497088 4012
rect 498256 3754 498284 4012
rect 499360 3754 499388 4012
rect 492460 3726 492536 3754
rect 493564 3726 493640 3754
rect 494760 3726 494836 3754
rect 495956 3726 496032 3754
rect 497060 3726 497136 3754
rect 498256 3726 498332 3754
rect 490104 1352 490156 1358
rect 490104 1294 490156 1300
rect 490748 1284 490800 1290
rect 490748 1226 490800 1232
rect 489000 1148 489052 1154
rect 489000 1090 489052 1096
rect 489920 944 489972 950
rect 489920 886 489972 892
rect 489932 480 489960 886
rect 487590 354 487702 480
rect 487264 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 1226
rect 491220 1086 491248 3726
rect 492508 1290 492536 3726
rect 493508 2848 493560 2854
rect 493508 2790 493560 2796
rect 492496 1284 492548 1290
rect 492496 1226 492548 1232
rect 492312 1216 492364 1222
rect 492312 1158 492364 1164
rect 491208 1080 491260 1086
rect 491208 1022 491260 1028
rect 492324 480 492352 1158
rect 493520 480 493548 2790
rect 493612 1222 493640 3726
rect 493600 1216 493652 1222
rect 493600 1158 493652 1164
rect 494704 1148 494756 1154
rect 494704 1090 494756 1096
rect 494716 480 494744 1090
rect 494808 678 494836 3726
rect 495532 1352 495584 1358
rect 495532 1294 495584 1300
rect 494796 672 494848 678
rect 494796 614 494848 620
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495544 354 495572 1294
rect 496004 1018 496032 3726
rect 497108 1358 497136 3726
rect 497096 1352 497148 1358
rect 497096 1294 497148 1300
rect 498304 1290 498332 3726
rect 499224 3726 499388 3754
rect 500556 3754 500584 4012
rect 501752 3754 501780 4012
rect 502856 3754 502884 4012
rect 504052 3754 504080 4012
rect 505156 3754 505184 4012
rect 506352 3754 506380 4012
rect 507548 3754 507576 4012
rect 500556 3726 500632 3754
rect 501752 3726 501828 3754
rect 502856 3726 502932 3754
rect 504052 3726 504128 3754
rect 505156 3726 505232 3754
rect 498200 1284 498252 1290
rect 498200 1226 498252 1232
rect 498292 1284 498344 1290
rect 498292 1226 498344 1232
rect 497096 1080 497148 1086
rect 497096 1022 497148 1028
rect 495992 1012 496044 1018
rect 495992 954 496044 960
rect 497108 480 497136 1022
rect 498212 480 498240 1226
rect 495870 354 495982 480
rect 495544 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499224 66 499252 3726
rect 500604 1222 500632 3726
rect 499396 1216 499448 1222
rect 499396 1158 499448 1164
rect 500592 1216 500644 1222
rect 500592 1158 500644 1164
rect 499408 480 499436 1158
rect 501800 1154 501828 3726
rect 501788 1148 501840 1154
rect 501788 1090 501840 1096
rect 502904 1018 502932 3726
rect 504100 1358 504128 3726
rect 502984 1352 503036 1358
rect 502984 1294 503036 1300
rect 504088 1352 504140 1358
rect 504088 1294 504140 1300
rect 501788 1012 501840 1018
rect 501788 954 501840 960
rect 502892 1012 502944 1018
rect 502892 954 502944 960
rect 500592 672 500644 678
rect 500592 614 500644 620
rect 500604 480 500632 614
rect 501800 480 501828 954
rect 502996 480 503024 1294
rect 503812 1284 503864 1290
rect 503812 1226 503864 1232
rect 499212 60 499264 66
rect 499212 2 499264 8
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503824 354 503852 1226
rect 505204 1086 505232 3726
rect 506308 3726 506380 3754
rect 507504 3726 507576 3754
rect 508652 3754 508680 4012
rect 509848 3754 509876 4012
rect 510952 3754 510980 4012
rect 512148 3754 512176 4012
rect 513344 3754 513372 4012
rect 508652 3726 508728 3754
rect 509848 3726 509924 3754
rect 510952 3726 511028 3754
rect 512148 3726 512224 3754
rect 505192 1080 505244 1086
rect 505192 1022 505244 1028
rect 504150 354 504262 480
rect 503824 326 504262 354
rect 504150 -960 504262 326
rect 505346 82 505458 480
rect 505346 66 505600 82
rect 506308 66 506336 3726
rect 506480 1216 506532 1222
rect 506480 1158 506532 1164
rect 506492 480 506520 1158
rect 507308 1148 507360 1154
rect 507308 1090 507360 1096
rect 505346 60 505612 66
rect 505346 54 505560 60
rect 505346 -960 505458 54
rect 505560 2 505612 8
rect 506296 60 506348 66
rect 506296 2 506348 8
rect 506450 -960 506562 480
rect 507320 82 507348 1090
rect 507504 202 507532 3726
rect 507492 196 507544 202
rect 507492 138 507544 144
rect 507646 82 507758 480
rect 508700 270 508728 3726
rect 509896 1358 509924 3726
rect 509700 1352 509752 1358
rect 509700 1294 509752 1300
rect 509884 1352 509936 1358
rect 509884 1294 509936 1300
rect 508872 1012 508924 1018
rect 508872 954 508924 960
rect 508884 480 508912 954
rect 508688 264 508740 270
rect 508688 206 508740 212
rect 507320 54 507758 82
rect 507646 -960 507758 54
rect 508842 -960 508954 480
rect 509712 354 509740 1294
rect 511000 1290 511028 3726
rect 510988 1284 511040 1290
rect 510988 1226 511040 1232
rect 512196 1086 512224 3726
rect 513300 3726 513372 3754
rect 514448 3754 514476 4012
rect 515644 3754 515672 4012
rect 516748 3754 516776 4012
rect 517944 3754 517972 4012
rect 519140 3754 519168 4012
rect 520244 3754 520272 4012
rect 514448 3726 514524 3754
rect 515644 3726 515720 3754
rect 516748 3726 516824 3754
rect 517944 3726 518020 3754
rect 519140 3726 519216 3754
rect 513300 1154 513328 3726
rect 513288 1148 513340 1154
rect 513288 1090 513340 1096
rect 511264 1080 511316 1086
rect 511264 1022 511316 1028
rect 512184 1080 512236 1086
rect 512184 1022 512236 1028
rect 511276 480 511304 1022
rect 514496 882 514524 3726
rect 514484 876 514536 882
rect 514484 818 514536 824
rect 510038 354 510150 480
rect 509712 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 82 512542 480
rect 513534 218 513646 480
rect 513392 202 513646 218
rect 513380 196 513646 202
rect 513432 190 513646 196
rect 513380 138 513432 144
rect 512104 66 512542 82
rect 512092 60 512542 66
rect 512144 54 512542 60
rect 512092 2 512144 8
rect 512430 -960 512542 54
rect 513534 -960 513646 190
rect 514730 218 514842 480
rect 514944 264 514996 270
rect 514730 212 514944 218
rect 514730 206 514996 212
rect 514730 190 514984 206
rect 514730 -960 514842 190
rect 515692 134 515720 3726
rect 515772 1352 515824 1358
rect 515772 1294 515824 1300
rect 515784 354 515812 1294
rect 515926 354 516038 480
rect 515784 326 516038 354
rect 515680 128 515732 134
rect 515680 70 515732 76
rect 515926 -960 516038 326
rect 516796 270 516824 3726
rect 517992 1290 518020 3726
rect 519188 1358 519216 3726
rect 520200 3726 520272 3754
rect 521440 3754 521468 4012
rect 522636 3754 522664 4012
rect 523740 3754 523768 4012
rect 524936 3754 524964 4012
rect 526040 3754 526068 4012
rect 527236 3754 527264 4012
rect 528432 3754 528460 4012
rect 529536 3754 529564 4012
rect 530732 3754 530760 4012
rect 531836 3754 531864 4012
rect 533032 3754 533060 4012
rect 534228 3754 534256 4012
rect 535332 3754 535360 4012
rect 536528 3754 536556 4012
rect 537632 3754 537660 4012
rect 538828 3754 538856 4012
rect 540024 3754 540052 4012
rect 541128 3754 541156 4012
rect 542324 3754 542352 4012
rect 521440 3726 521516 3754
rect 522636 3726 522712 3754
rect 523740 3726 523816 3754
rect 524936 3726 525012 3754
rect 526040 3726 526116 3754
rect 527236 3726 527312 3754
rect 528432 3726 528508 3754
rect 529536 3726 529612 3754
rect 530732 3726 530808 3754
rect 531836 3726 531912 3754
rect 533032 3726 533108 3754
rect 534228 3726 534304 3754
rect 535332 3726 535408 3754
rect 536528 3726 536604 3754
rect 537632 3726 537708 3754
rect 538828 3726 538904 3754
rect 540024 3726 540100 3754
rect 541128 3726 541204 3754
rect 519176 1352 519228 1358
rect 519176 1294 519228 1300
rect 517152 1284 517204 1290
rect 517152 1226 517204 1232
rect 517980 1284 518032 1290
rect 517980 1226 518032 1232
rect 517164 480 517192 1226
rect 519544 1148 519596 1154
rect 519544 1090 519596 1096
rect 517980 1080 518032 1086
rect 517980 1022 518032 1028
rect 516784 264 516836 270
rect 516784 206 516836 212
rect 517122 -960 517234 480
rect 517992 354 518020 1022
rect 519556 480 519584 1090
rect 520200 1086 520228 3726
rect 520188 1080 520240 1086
rect 520188 1022 520240 1028
rect 521488 882 521516 3726
rect 522684 1222 522712 3726
rect 522672 1216 522724 1222
rect 522672 1158 522724 1164
rect 523788 1154 523816 3726
rect 523868 1284 523920 1290
rect 523868 1226 523920 1232
rect 523776 1148 523828 1154
rect 523776 1090 523828 1096
rect 520740 876 520792 882
rect 520740 818 520792 824
rect 521476 876 521528 882
rect 521476 818 521528 824
rect 520752 480 520780 818
rect 518318 354 518430 480
rect 517992 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521660 128 521712 134
rect 521814 82 521926 480
rect 521712 76 521926 82
rect 521660 70 521926 76
rect 521672 54 521926 70
rect 521814 -960 521926 54
rect 523010 218 523122 480
rect 523880 354 523908 1226
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 523224 264 523276 270
rect 523010 212 523224 218
rect 523010 206 523276 212
rect 523010 190 523264 206
rect 523010 -960 523122 190
rect 524206 -960 524318 326
rect 524984 134 525012 3726
rect 526088 1358 526116 3726
rect 525432 1352 525484 1358
rect 525432 1294 525484 1300
rect 526076 1352 526128 1358
rect 526076 1294 526128 1300
rect 525444 480 525472 1294
rect 527284 1290 527312 3726
rect 527272 1284 527324 1290
rect 527272 1226 527324 1232
rect 526628 1080 526680 1086
rect 526628 1022 526680 1028
rect 526640 480 526668 1022
rect 527824 876 527876 882
rect 527824 818 527876 824
rect 527836 480 527864 818
rect 524972 128 525024 134
rect 524972 70 525024 76
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528480 66 528508 3726
rect 529020 1216 529072 1222
rect 529020 1158 529072 1164
rect 529032 480 529060 1158
rect 529584 1086 529612 3726
rect 530780 1222 530808 3726
rect 530768 1216 530820 1222
rect 530768 1158 530820 1164
rect 530124 1148 530176 1154
rect 530124 1090 530176 1096
rect 529572 1080 529624 1086
rect 529572 1022 529624 1028
rect 530136 480 530164 1090
rect 531884 610 531912 3726
rect 532148 1352 532200 1358
rect 532148 1294 532200 1300
rect 531872 604 531924 610
rect 531872 546 531924 552
rect 528468 60 528520 66
rect 528468 2 528520 8
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 82 531402 480
rect 532160 354 532188 1294
rect 533080 1154 533108 3726
rect 534276 1358 534304 3726
rect 534264 1352 534316 1358
rect 534264 1294 534316 1300
rect 533712 1284 533764 1290
rect 533712 1226 533764 1232
rect 533068 1148 533120 1154
rect 533068 1090 533120 1096
rect 533724 480 533752 1226
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 531504 128 531556 134
rect 531290 76 531504 82
rect 531290 70 531556 76
rect 531290 54 531544 70
rect 531290 -960 531402 54
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534878 82 534990 480
rect 535380 474 535408 3726
rect 536104 1080 536156 1086
rect 536104 1022 536156 1028
rect 536116 480 536144 1022
rect 535368 468 535420 474
rect 535368 410 535420 416
rect 534552 66 534990 82
rect 534540 60 534990 66
rect 534592 54 534990 60
rect 534540 2 534592 8
rect 534878 -960 534990 54
rect 536074 -960 536186 480
rect 536576 66 536604 3726
rect 537208 1216 537260 1222
rect 537208 1158 537260 1164
rect 537220 480 537248 1158
rect 537680 542 537708 3726
rect 538876 1222 538904 3726
rect 538864 1216 538916 1222
rect 538864 1158 538916 1164
rect 539600 1148 539652 1154
rect 539600 1090 539652 1096
rect 538404 604 538456 610
rect 538404 546 538456 552
rect 537668 536 537720 542
rect 536564 60 536616 66
rect 536564 2 536616 8
rect 537178 -960 537290 480
rect 537668 478 537720 484
rect 538416 480 538444 546
rect 539612 480 539640 1090
rect 540072 1018 540100 3726
rect 540428 1352 540480 1358
rect 540428 1294 540480 1300
rect 540060 1012 540112 1018
rect 540060 954 540112 960
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540440 354 540468 1294
rect 541176 1290 541204 3726
rect 542280 3726 542352 3754
rect 543428 3754 543456 4012
rect 544624 3754 544652 4012
rect 545820 3754 545848 4012
rect 546924 3754 546952 4012
rect 548120 3754 548148 4012
rect 549316 3754 549344 4012
rect 550420 3754 550448 4012
rect 551616 3754 551644 4012
rect 552720 3754 552748 4012
rect 553916 3754 553944 4012
rect 555112 3754 555140 4012
rect 556216 3754 556244 4012
rect 557412 3754 557440 4012
rect 558516 3754 558544 4012
rect 559712 3754 559740 4012
rect 543428 3726 543504 3754
rect 544624 3726 544700 3754
rect 545820 3726 545896 3754
rect 546924 3726 547000 3754
rect 548120 3726 548196 3754
rect 549316 3726 549392 3754
rect 550420 3726 550496 3754
rect 551616 3726 551692 3754
rect 552720 3726 552796 3754
rect 553916 3726 553992 3754
rect 555112 3726 555188 3754
rect 556216 3726 556292 3754
rect 557412 3726 557488 3754
rect 542280 1358 542308 3726
rect 542268 1352 542320 1358
rect 542268 1294 542320 1300
rect 541164 1284 541216 1290
rect 541164 1226 541216 1232
rect 543476 1154 543504 3726
rect 543464 1148 543516 1154
rect 543464 1090 543516 1096
rect 544672 746 544700 3726
rect 545488 1216 545540 1222
rect 545488 1158 545540 1164
rect 544660 740 544712 746
rect 544660 682 544712 688
rect 544384 604 544436 610
rect 544384 546 544436 552
rect 544396 480 544424 546
rect 545500 480 545528 1158
rect 545868 1086 545896 3726
rect 545856 1080 545908 1086
rect 545856 1022 545908 1028
rect 546684 1012 546736 1018
rect 546684 954 546736 960
rect 546696 480 546724 954
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 354 542074 480
rect 542176 468 542228 474
rect 542176 410 542228 416
rect 542188 354 542216 410
rect 541962 326 542216 354
rect 541962 -960 542074 326
rect 543158 82 543270 480
rect 542832 66 543270 82
rect 542820 60 543270 66
rect 542872 54 543270 60
rect 542820 2 542872 8
rect 543158 -960 543270 54
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 546972 66 547000 3726
rect 548168 1290 548196 3726
rect 549076 1352 549128 1358
rect 549076 1294 549128 1300
rect 547880 1284 547932 1290
rect 547880 1226 547932 1232
rect 548156 1284 548208 1290
rect 548156 1226 548208 1232
rect 547892 480 547920 1226
rect 549088 480 549116 1294
rect 549364 610 549392 3726
rect 550468 1222 550496 3726
rect 551664 1358 551692 3726
rect 551652 1352 551704 1358
rect 551652 1294 551704 1300
rect 550456 1216 550508 1222
rect 550456 1158 550508 1164
rect 552768 1154 552796 3726
rect 550272 1148 550324 1154
rect 550272 1090 550324 1096
rect 552756 1148 552808 1154
rect 552756 1090 552808 1096
rect 549352 604 549404 610
rect 549352 546 549404 552
rect 550284 480 550312 1090
rect 552664 1080 552716 1086
rect 552664 1022 552716 1028
rect 551468 740 551520 746
rect 551468 682 551520 688
rect 551480 480 551508 682
rect 552676 480 552704 1022
rect 546960 60 547012 66
rect 546960 2 547012 8
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 82 553850 480
rect 553964 270 553992 3726
rect 554964 1284 555016 1290
rect 554964 1226 555016 1232
rect 554976 480 555004 1226
rect 555160 746 555188 3726
rect 555148 740 555200 746
rect 555148 682 555200 688
rect 556264 678 556292 3726
rect 557356 1216 557408 1222
rect 557356 1158 557408 1164
rect 556252 672 556304 678
rect 556252 614 556304 620
rect 556160 604 556212 610
rect 556160 546 556212 552
rect 556172 480 556200 546
rect 557368 480 557396 1158
rect 557460 626 557488 3726
rect 558472 3726 558544 3754
rect 559668 3726 559740 3754
rect 560908 3754 560936 4012
rect 562012 3754 562040 4012
rect 563208 3754 563236 4012
rect 564312 3754 564340 4012
rect 565508 3754 565536 4012
rect 566704 3754 566732 4012
rect 560908 3726 560984 3754
rect 562012 3726 562088 3754
rect 563208 3726 563376 3754
rect 558472 1222 558500 3726
rect 558552 1352 558604 1358
rect 558552 1294 558604 1300
rect 558460 1216 558512 1222
rect 558460 1158 558512 1164
rect 557460 598 557580 626
rect 557552 542 557580 598
rect 557540 536 557592 542
rect 553952 264 554004 270
rect 553952 206 554004 212
rect 553738 66 553992 82
rect 553738 60 554004 66
rect 553738 54 553952 60
rect 553738 -960 553850 54
rect 553952 2 554004 8
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 557540 478 557592 484
rect 558564 480 558592 1294
rect 559668 1086 559696 3726
rect 560956 1358 560984 3726
rect 560944 1352 560996 1358
rect 560944 1294 560996 1300
rect 562060 1290 562088 3726
rect 562048 1284 562100 1290
rect 562048 1226 562100 1232
rect 559748 1148 559800 1154
rect 559748 1090 559800 1096
rect 559656 1080 559708 1086
rect 559656 1022 559708 1028
rect 559760 480 559788 1090
rect 562048 740 562100 746
rect 562048 682 562100 688
rect 562060 480 562088 682
rect 563152 672 563204 678
rect 563204 620 563284 626
rect 563152 614 563284 620
rect 563164 598 563284 614
rect 563348 610 563376 3726
rect 564268 3726 564340 3754
rect 565464 3726 565536 3754
rect 566660 3726 566732 3754
rect 567808 3754 567836 4012
rect 569004 3754 569032 4012
rect 570108 3754 570136 4012
rect 571304 3754 571332 4012
rect 567808 3726 567884 3754
rect 569004 3726 569080 3754
rect 570108 3726 570184 3754
rect 563256 480 563284 598
rect 563336 604 563388 610
rect 563336 546 563388 552
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560484 264 560536 270
rect 560822 218 560934 480
rect 560536 212 560934 218
rect 560484 206 560934 212
rect 560496 190 560934 206
rect 560822 -960 560934 190
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564268 270 564296 3726
rect 564624 536 564676 542
rect 564410 354 564522 480
rect 564624 478 564676 484
rect 564636 354 564664 478
rect 564410 326 564664 354
rect 565464 338 565492 3726
rect 565636 1216 565688 1222
rect 565636 1158 565688 1164
rect 565648 480 565676 1158
rect 565452 332 565504 338
rect 564256 264 564308 270
rect 564256 206 564308 212
rect 564410 -960 564522 326
rect 565452 274 565504 280
rect 565606 -960 565718 480
rect 566660 474 566688 3726
rect 567856 1154 567884 3726
rect 568028 1352 568080 1358
rect 568028 1294 568080 1300
rect 567844 1148 567896 1154
rect 567844 1090 567896 1096
rect 566832 1080 566884 1086
rect 566832 1022 566884 1028
rect 566844 480 566872 1022
rect 568040 480 568068 1294
rect 569052 1222 569080 3726
rect 570156 1290 570184 3726
rect 571260 3726 571332 3754
rect 572500 3754 572528 4012
rect 573604 3754 573632 4012
rect 574800 3754 574828 4012
rect 575918 3998 576164 4026
rect 572500 3726 572576 3754
rect 573604 3726 573680 3754
rect 574800 3726 574876 3754
rect 571260 1358 571288 3726
rect 571248 1352 571300 1358
rect 571248 1294 571300 1300
rect 569132 1284 569184 1290
rect 569132 1226 569184 1232
rect 570144 1284 570196 1290
rect 570144 1226 570196 1232
rect 569040 1216 569092 1222
rect 569040 1158 569092 1164
rect 569144 480 569172 1226
rect 570328 604 570380 610
rect 570328 546 570380 552
rect 570340 480 570368 546
rect 566648 468 566700 474
rect 566648 410 566700 416
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571340 264 571392 270
rect 571494 218 571606 480
rect 571392 212 571606 218
rect 571340 206 571606 212
rect 571352 190 571606 206
rect 571494 -960 571606 190
rect 572548 66 572576 3726
rect 572690 354 572802 480
rect 572690 338 572944 354
rect 572690 332 572956 338
rect 572690 326 572904 332
rect 572536 60 572588 66
rect 572536 2 572588 8
rect 572690 -960 572802 326
rect 572904 274 572956 280
rect 573652 134 573680 3726
rect 573732 468 573784 474
rect 573732 410 573784 416
rect 573744 354 573772 410
rect 573886 354 573998 480
rect 573744 326 573998 354
rect 573640 128 573692 134
rect 573640 70 573692 76
rect 573886 -960 573998 326
rect 574848 270 574876 3726
rect 575112 1148 575164 1154
rect 575112 1090 575164 1096
rect 575124 480 575152 1090
rect 574836 264 574888 270
rect 574836 206 574888 212
rect 575082 -960 575194 480
rect 576136 338 576164 3998
rect 578608 1352 578660 1358
rect 578608 1294 578660 1300
rect 577412 1284 577464 1290
rect 577412 1226 577464 1232
rect 576308 1216 576360 1222
rect 576308 1158 576360 1164
rect 576320 480 576348 1158
rect 577424 480 577452 1226
rect 578620 480 578648 1294
rect 576124 332 576176 338
rect 576124 274 576176 280
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 82 579886 480
rect 579632 66 579886 82
rect 579620 60 579886 66
rect 579672 54 579886 60
rect 579620 2 579672 8
rect 579774 -960 579886 54
rect 580970 82 581082 480
rect 581828 264 581880 270
rect 582166 218 582278 480
rect 581880 212 582278 218
rect 581828 206 582278 212
rect 581840 190 582278 206
rect 581184 128 581236 134
rect 580970 76 581184 82
rect 580970 70 581236 76
rect 580970 54 581224 70
rect 580970 -960 581082 54
rect 582166 -960 582278 190
rect 583362 354 583474 480
rect 583362 338 583616 354
rect 583362 332 583628 338
rect 583362 326 583576 332
rect 583362 -960 583474 326
rect 583576 274 583628 280
<< via2 >>
rect 3514 697920 3570 697976
rect 3514 697312 3570 697368
rect 579526 684664 579582 684720
rect 579618 683848 579674 683904
rect 578330 644564 578386 644600
rect 578330 644544 578332 644564
rect 578332 644544 578384 644564
rect 578384 644544 578386 644564
rect 580906 644000 580962 644056
rect 3422 436600 3478 436656
rect 3422 435986 3478 436042
rect 3422 423544 3478 423600
rect 3422 422932 3478 422988
rect 3422 410488 3478 410544
rect 3422 409878 3478 409934
rect 3422 397432 3478 397488
rect 3422 396824 3478 396880
rect 3422 384376 3478 384432
rect 3422 383648 3478 383704
rect 3422 371320 3478 371376
rect 3422 370594 3478 370650
rect 3422 358400 3478 358456
rect 3422 357540 3478 357596
rect 579526 351872 579582 351928
rect 579526 351056 579582 351112
rect 3422 345344 3478 345400
rect 3422 344364 3478 344420
rect 579618 338544 579674 338600
rect 579526 337864 579582 337920
rect 3422 332288 3478 332344
rect 3422 331310 3478 331366
rect 580170 325216 580226 325272
rect 580170 324400 580226 324456
rect 3422 319232 3478 319288
rect 3422 318256 3478 318312
rect 579618 312024 579674 312080
rect 579526 311072 579582 311128
rect 3422 306176 3478 306232
rect 3422 305080 3478 305136
rect 579618 298696 579674 298752
rect 579526 297744 579582 297800
rect 3422 293120 3478 293176
rect 3422 292026 3478 292082
rect 580170 285368 580226 285424
rect 580170 284416 580226 284472
rect 3422 280064 3478 280120
rect 3422 278972 3478 279028
rect 579618 272176 579674 272232
rect 579526 271088 579582 271144
rect 3422 267144 3478 267200
rect 3422 265918 3478 265974
rect 580906 258848 580962 258904
rect 578882 257624 578938 257680
rect 3422 254088 3478 254144
rect 3422 252742 3478 252798
rect 580170 245520 580226 245576
rect 580170 244432 580226 244488
rect 3422 241032 3478 241088
rect 3422 239688 3478 239744
rect 579618 232328 579674 232384
rect 579526 231104 579582 231160
rect 3422 227976 3478 228032
rect 3422 226634 3478 226690
rect 579618 219000 579674 219056
rect 579526 217640 579582 217696
rect 3422 214920 3478 214976
rect 3422 213458 3478 213514
rect 579618 205672 579674 205728
rect 579526 204312 579582 204368
rect 3422 201864 3478 201920
rect 3422 200404 3478 200460
rect 579618 192480 579674 192536
rect 579526 190984 579582 191040
rect 3606 188808 3662 188864
rect 3606 187350 3662 187406
rect 579618 179152 579674 179208
rect 579526 177656 579582 177712
rect 3422 175888 3478 175944
rect 3422 174174 3478 174230
rect 579618 165824 579674 165880
rect 579526 164328 579582 164384
rect 2134 162832 2190 162888
rect 2134 161064 2190 161120
rect 580906 152632 580962 152688
rect 578514 151000 578570 151056
rect 3422 149776 3478 149832
rect 3422 148066 3478 148122
rect 579618 139304 579674 139360
rect 579526 137536 579582 137592
rect 2134 136720 2190 136776
rect 2134 134952 2190 135008
rect 579618 125976 579674 126032
rect 579526 124344 579582 124400
rect 3422 123664 3478 123720
rect 3422 121836 3478 121892
rect 579618 112784 579674 112840
rect 579526 110880 579582 110936
rect 2134 110608 2190 110664
rect 2134 108840 2190 108896
rect 579618 99456 579674 99512
rect 3422 97552 3478 97608
rect 579526 97552 579582 97608
rect 3422 95728 3478 95784
rect 579618 86128 579674 86184
rect 2134 84632 2190 84688
rect 579526 84224 579582 84280
rect 2134 82592 2190 82648
rect 579618 72936 579674 72992
rect 3422 71576 3478 71632
rect 579526 70896 579582 70952
rect 3422 69498 3478 69554
rect 579618 59608 579674 59664
rect 2134 58520 2190 58576
rect 579526 57568 579582 57624
rect 2134 56480 2190 56536
rect 579986 46280 580042 46336
rect 3422 45464 3478 45520
rect 578330 44240 578386 44296
rect 3422 43268 3478 43324
rect 579618 33088 579674 33144
rect 2134 32408 2190 32464
rect 579526 30912 579582 30968
rect 2134 30232 2190 30288
rect 579618 19760 579674 19816
rect 2042 19352 2098 19408
rect 579526 17584 579582 17640
rect 2042 17176 2098 17232
rect 579618 6568 579674 6624
rect 2778 6432 2834 6488
rect 2778 4120 2834 4176
rect 579526 4120 579582 4176
<< metal3 >>
rect 3509 697978 3575 697981
rect 3509 697976 4048 697978
rect 3509 697920 3514 697976
rect 3570 697920 4048 697976
rect 3509 697918 4048 697920
rect 575920 697918 576410 697978
rect 3509 697915 3575 697918
rect 576350 697914 576410 697918
rect 576350 697854 583586 697914
rect -960 697370 480 697460
rect 3509 697370 3575 697373
rect 583526 697370 583586 697854
rect -960 697368 3575 697370
rect -960 697312 3514 697368
rect 3570 697312 3575 697368
rect -960 697310 3575 697312
rect -960 697220 480 697310
rect 3509 697307 3575 697310
rect 583342 697324 583586 697370
rect 583342 697310 584960 697324
rect 583342 697234 583402 697310
rect 583520 697234 584960 697310
rect 583342 697174 584960 697234
rect 583520 697084 584960 697174
rect 3374 684742 4048 684802
rect -960 684314 480 684404
rect 3374 684314 3434 684742
rect 579521 684722 579587 684725
rect 576350 684720 579587 684722
rect 576350 684680 579526 684720
rect 575920 684664 579526 684680
rect 579582 684664 579587 684720
rect 575920 684662 579587 684664
rect 575920 684620 576410 684662
rect 579521 684659 579587 684662
rect -960 684254 3434 684314
rect -960 684164 480 684254
rect 579613 683906 579679 683909
rect 583520 683906 584960 683996
rect 579613 683904 584960 683906
rect 579613 683848 579618 683904
rect 579674 683848 584960 683904
rect 579613 683846 584960 683848
rect 579613 683843 579679 683846
rect 583520 683756 584960 683846
rect 3374 671688 4048 671748
rect -960 671258 480 671348
rect 3374 671258 3434 671688
rect 576350 671382 583586 671394
rect 575920 671334 583586 671382
rect 575920 671322 576410 671334
rect -960 671198 3434 671258
rect -960 671108 480 671198
rect 583526 670850 583586 671334
rect 583342 670804 583586 670850
rect 583342 670790 584960 670804
rect 583342 670714 583402 670790
rect 583520 670714 584960 670790
rect 583342 670654 584960 670714
rect 583520 670564 584960 670654
rect 3374 658634 4048 658694
rect -960 658202 480 658292
rect 3374 658202 3434 658634
rect -960 658142 3434 658202
rect -960 658052 480 658142
rect 575920 657930 576410 657962
rect 575920 657902 583586 657930
rect 576350 657870 583586 657902
rect 583526 657522 583586 657870
rect 583342 657476 583586 657522
rect 583342 657462 584960 657476
rect 583342 657386 583402 657462
rect 583520 657386 584960 657462
rect 583342 657326 584960 657386
rect 583520 657236 584960 657326
rect 3374 645458 4048 645518
rect -960 645146 480 645236
rect 3374 645146 3434 645458
rect -960 645086 3434 645146
rect -960 644996 480 645086
rect 575920 644604 576410 644664
rect 576350 644602 576410 644604
rect 578325 644602 578391 644605
rect 576350 644600 578391 644602
rect 576350 644544 578330 644600
rect 578386 644544 578391 644600
rect 576350 644542 578391 644544
rect 578325 644539 578391 644542
rect 580901 644058 580967 644061
rect 583520 644058 584960 644148
rect 580901 644056 584960 644058
rect 580901 644000 580906 644056
rect 580962 644000 584960 644056
rect 580901 643998 584960 644000
rect 580901 643995 580967 643998
rect 583520 643908 584960 643998
rect 3374 632404 4048 632464
rect -960 632090 480 632180
rect 3374 632090 3434 632404
rect -960 632030 3434 632090
rect -960 631940 480 632030
rect 575920 631306 576410 631366
rect 576350 631274 576410 631306
rect 576350 631214 583586 631274
rect 583526 631002 583586 631214
rect 583342 630956 583586 631002
rect 583342 630942 584960 630956
rect 583342 630866 583402 630942
rect 583520 630866 584960 630942
rect 583342 630806 584960 630866
rect 583520 630716 584960 630806
rect 3374 619350 4048 619410
rect -960 619170 480 619260
rect 3374 619170 3434 619350
rect -960 619110 3434 619170
rect -960 619020 480 619110
rect 575920 617886 583586 617946
rect 583526 617674 583586 617886
rect 583342 617628 583586 617674
rect 583342 617614 584960 617628
rect 583342 617538 583402 617614
rect 583520 617538 584960 617614
rect 583342 617478 584960 617538
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3374 606174 4048 606234
rect 3374 606114 3434 606174
rect -960 606054 3434 606114
rect -960 605964 480 606054
rect 575920 604618 576410 604648
rect 575920 604588 576870 604618
rect 576350 604558 576870 604588
rect 576810 604482 576870 604558
rect 576810 604422 579722 604482
rect 579662 604210 579722 604422
rect 583520 604210 584960 604300
rect 579662 604150 584960 604210
rect 583520 604060 584960 604150
rect -960 593058 480 593148
rect 3374 593120 4048 593180
rect 3374 593058 3434 593120
rect -960 592998 3434 593058
rect -960 592908 480 592998
rect 575920 591290 576410 591350
rect 576350 591230 576870 591290
rect 576810 591018 576870 591230
rect 583520 591018 584960 591108
rect 576810 590958 584960 591018
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3374 580066 4048 580126
rect 3374 580002 3434 580066
rect -960 579942 3434 580002
rect -960 579852 480 579942
rect 575920 577870 576410 577930
rect 576350 577826 576410 577870
rect 576350 577766 576870 577826
rect 576810 577690 576870 577766
rect 583520 577690 584960 577780
rect 576810 577630 584960 577690
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3374 566946 4048 566950
rect -960 566890 4048 566946
rect -960 566886 3434 566890
rect -960 566796 480 566886
rect 575920 564572 576410 564632
rect 576350 564498 576410 564572
rect 576350 564438 579722 564498
rect 579662 564362 579722 564438
rect 583520 564362 584960 564452
rect 579662 564302 584960 564362
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3374 553890 4048 553896
rect -960 553836 4048 553890
rect -960 553830 3434 553836
rect -960 553740 480 553830
rect 575920 551170 576410 551212
rect 583520 551170 584960 551260
rect 575920 551152 584960 551170
rect 576350 551110 584960 551152
rect 583520 551020 584960 551110
rect -960 540834 480 540924
rect 3374 540834 4048 540842
rect -960 540782 4048 540834
rect -960 540774 3434 540782
rect -960 540684 480 540774
rect 575920 537854 576410 537914
rect 576350 537842 576410 537854
rect 583520 537842 584960 537932
rect 576350 537782 584960 537842
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect -960 527854 3434 527914
rect -960 527764 480 527854
rect 3374 527788 3434 527854
rect 3374 527728 4048 527788
rect 575920 524556 576410 524616
rect 576350 524514 576410 524556
rect 583520 524514 584960 524604
rect 576350 524454 584960 524514
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect -960 514798 3434 514858
rect -960 514708 480 514798
rect 3374 514612 3434 514798
rect 3374 514552 4048 514612
rect 583520 511322 584960 511412
rect 576350 511262 584960 511322
rect 576350 511196 576410 511262
rect 575920 511136 576410 511196
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect -960 501742 3434 501802
rect -960 501652 480 501742
rect 3374 501558 3434 501742
rect 3374 501498 4048 501558
rect 583520 497994 584960 498084
rect 576350 497934 584960 497994
rect 576350 497898 576410 497934
rect 575920 497838 576410 497898
rect 583520 497844 584960 497934
rect -960 488746 480 488836
rect -960 488686 3434 488746
rect -960 488596 480 488686
rect 3374 488504 3434 488686
rect 3374 488444 4048 488504
rect 583520 484666 584960 484756
rect 576350 484606 584960 484666
rect 576350 484600 576410 484606
rect 575920 484540 576410 484600
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect -960 475630 3434 475690
rect -960 475540 480 475630
rect 3374 475328 3434 475630
rect 3374 475268 4048 475328
rect 583520 471474 584960 471564
rect 576810 471414 584960 471474
rect 576810 471202 576870 471414
rect 583520 471324 584960 471414
rect 576350 471180 576870 471202
rect 575920 471142 576870 471180
rect 575920 471120 576410 471142
rect -960 462634 480 462724
rect -960 462574 3434 462634
rect -960 462484 480 462574
rect 3374 462274 3434 462574
rect 3374 462214 4048 462274
rect 583520 458146 584960 458236
rect 576810 458086 584960 458146
rect 576810 458010 576870 458086
rect 576350 457950 576870 458010
rect 583520 457996 584960 458086
rect 576350 457882 576410 457950
rect 575920 457822 576410 457882
rect -960 449578 480 449668
rect -960 449518 3434 449578
rect -960 449428 480 449518
rect 3374 449220 3434 449518
rect 3374 449160 4048 449220
rect 583520 444818 584960 444908
rect 576810 444758 584960 444818
rect 576810 444682 576870 444758
rect 576350 444622 576870 444682
rect 583520 444668 584960 444758
rect 576350 444584 576410 444622
rect 575920 444524 576410 444584
rect -960 436658 480 436748
rect 3417 436658 3483 436661
rect -960 436656 3483 436658
rect -960 436600 3422 436656
rect 3478 436600 3483 436656
rect -960 436598 3483 436600
rect -960 436508 480 436598
rect 3417 436595 3483 436598
rect 3417 436044 3483 436047
rect 3417 436042 4048 436044
rect 3417 435986 3422 436042
rect 3478 435986 4048 436042
rect 3417 435984 4048 435986
rect 3417 435981 3483 435984
rect 583520 431626 584960 431716
rect 583342 431566 584960 431626
rect 583342 431490 583402 431566
rect 583520 431490 584960 431566
rect 583342 431476 584960 431490
rect 583342 431430 583586 431476
rect 583526 431218 583586 431430
rect 576350 431164 583586 431218
rect 575920 431158 583586 431164
rect 575920 431104 576410 431158
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 3417 422990 3483 422993
rect 3417 422988 4048 422990
rect 3417 422932 3422 422988
rect 3478 422932 4048 422988
rect 3417 422930 4048 422932
rect 3417 422927 3483 422930
rect 583520 418298 584960 418388
rect 579662 418238 584960 418298
rect 579662 418162 579722 418238
rect 576810 418102 579722 418162
rect 583520 418148 584960 418238
rect 576810 417890 576870 418102
rect 576350 417866 576870 417890
rect 575920 417830 576870 417866
rect 575920 417806 576410 417830
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 3417 409936 3483 409939
rect 3417 409934 4048 409936
rect 3417 409878 3422 409934
rect 3478 409878 4048 409934
rect 3417 409876 4048 409878
rect 3417 409873 3483 409876
rect 583520 404970 584960 405060
rect 583342 404910 584960 404970
rect 583342 404834 583402 404910
rect 583520 404834 584960 404910
rect 583342 404820 584960 404834
rect 583342 404774 583586 404820
rect 583526 404562 583586 404774
rect 576350 404502 583586 404562
rect 576350 404446 576410 404502
rect 575920 404386 576410 404446
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 3417 396882 3483 396885
rect 3417 396880 4048 396882
rect 3417 396824 3422 396880
rect 3478 396824 4048 396880
rect 3417 396822 4048 396824
rect 3417 396819 3483 396822
rect 583520 391778 584960 391868
rect 583342 391718 584960 391778
rect 583342 391642 583402 391718
rect 583520 391642 584960 391718
rect 583342 391628 584960 391642
rect 583342 391582 583586 391628
rect 583526 391234 583586 391582
rect 576350 391174 583586 391234
rect 576350 391148 576410 391174
rect 575920 391088 576410 391148
rect -960 384434 480 384524
rect 3417 384434 3483 384437
rect -960 384432 3483 384434
rect -960 384376 3422 384432
rect 3478 384376 3483 384432
rect -960 384374 3483 384376
rect -960 384284 480 384374
rect 3417 384371 3483 384374
rect 3417 383706 3483 383709
rect 3417 383704 4048 383706
rect 3417 383648 3422 383704
rect 3478 383648 4048 383704
rect 3417 383646 4048 383648
rect 3417 383643 3483 383646
rect 583520 378450 584960 378540
rect 579662 378390 584960 378450
rect 579662 378178 579722 378390
rect 583520 378300 584960 378390
rect 579478 378118 579722 378178
rect 579478 377906 579538 378118
rect 576350 377850 579538 377906
rect 575920 377846 579538 377850
rect 575920 377790 576410 377846
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 3417 370652 3483 370655
rect 3417 370650 4048 370652
rect 3417 370594 3422 370650
rect 3478 370594 4048 370650
rect 3417 370592 4048 370594
rect 3417 370589 3483 370592
rect 583520 365122 584960 365212
rect 583342 365062 584960 365122
rect 583342 364986 583402 365062
rect 583520 364986 584960 365062
rect 583342 364972 584960 364986
rect 583342 364926 583586 364972
rect 583526 364442 583586 364926
rect 576350 364430 583586 364442
rect 575920 364382 583586 364430
rect 575920 364370 576410 364382
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 3417 357598 3483 357601
rect 3417 357596 4048 357598
rect 3417 357540 3422 357596
rect 3478 357540 4048 357596
rect 3417 357538 4048 357540
rect 3417 357535 3483 357538
rect 579521 351930 579587 351933
rect 583520 351930 584960 352020
rect 579521 351928 584960 351930
rect 579521 351872 579526 351928
rect 579582 351872 584960 351928
rect 579521 351870 584960 351872
rect 579521 351867 579587 351870
rect 583520 351780 584960 351870
rect 575920 351114 576410 351132
rect 579521 351114 579587 351117
rect 575920 351112 579587 351114
rect 575920 351072 579526 351112
rect 576350 351056 579526 351072
rect 579582 351056 579587 351112
rect 576350 351054 579587 351056
rect 579521 351051 579587 351054
rect -960 345402 480 345492
rect 3417 345402 3483 345405
rect -960 345400 3483 345402
rect -960 345344 3422 345400
rect 3478 345344 3483 345400
rect -960 345342 3483 345344
rect -960 345252 480 345342
rect 3417 345339 3483 345342
rect 3417 344422 3483 344425
rect 3417 344420 4048 344422
rect 3417 344364 3422 344420
rect 3478 344364 4048 344420
rect 3417 344362 4048 344364
rect 3417 344359 3483 344362
rect 579613 338602 579679 338605
rect 583520 338602 584960 338692
rect 579613 338600 584960 338602
rect 579613 338544 579618 338600
rect 579674 338544 584960 338600
rect 579613 338542 584960 338544
rect 579613 338539 579679 338542
rect 583520 338452 584960 338542
rect 579521 337922 579587 337925
rect 576350 337920 579587 337922
rect 576350 337864 579526 337920
rect 579582 337864 579587 337920
rect 576350 337862 579587 337864
rect 576350 337834 576410 337862
rect 579521 337859 579587 337862
rect 575920 337774 576410 337834
rect -960 332346 480 332436
rect 3417 332346 3483 332349
rect -960 332344 3483 332346
rect -960 332288 3422 332344
rect 3478 332288 3483 332344
rect -960 332286 3483 332288
rect -960 332196 480 332286
rect 3417 332283 3483 332286
rect 3417 331368 3483 331371
rect 3417 331366 4048 331368
rect 3417 331310 3422 331366
rect 3478 331310 4048 331366
rect 3417 331308 4048 331310
rect 3417 331305 3483 331308
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 580165 324458 580231 324461
rect 576350 324456 580231 324458
rect 576350 324414 580170 324456
rect 575920 324400 580170 324414
rect 580226 324400 580231 324456
rect 575920 324398 580231 324400
rect 575920 324354 576410 324398
rect 580165 324395 580231 324398
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 3417 318314 3483 318317
rect 3417 318312 4048 318314
rect 3417 318256 3422 318312
rect 3478 318256 4048 318312
rect 3417 318254 4048 318256
rect 3417 318251 3483 318254
rect 579613 312082 579679 312085
rect 583520 312082 584960 312172
rect 579613 312080 584960 312082
rect 579613 312024 579618 312080
rect 579674 312024 584960 312080
rect 579613 312022 584960 312024
rect 579613 312019 579679 312022
rect 583520 311932 584960 312022
rect 579521 311130 579587 311133
rect 576350 311128 579587 311130
rect 576350 311116 579526 311128
rect 575920 311072 579526 311116
rect 579582 311072 579587 311128
rect 575920 311070 579587 311072
rect 575920 311056 576410 311070
rect 579521 311067 579587 311070
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 3417 305138 3483 305141
rect 3417 305136 4048 305138
rect 3417 305080 3422 305136
rect 3478 305080 4048 305136
rect 3417 305078 4048 305080
rect 3417 305075 3483 305078
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect 575920 297802 576410 297818
rect 579521 297802 579587 297805
rect 575920 297800 579587 297802
rect 575920 297758 579526 297800
rect 576350 297744 579526 297758
rect 579582 297744 579587 297800
rect 576350 297742 579587 297744
rect 579521 297739 579587 297742
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 3417 292084 3483 292087
rect 3417 292082 4048 292084
rect 3417 292026 3422 292082
rect 3478 292026 4048 292082
rect 3417 292024 4048 292026
rect 3417 292021 3483 292024
rect 580165 285426 580231 285429
rect 583520 285426 584960 285516
rect 580165 285424 584960 285426
rect 580165 285368 580170 285424
rect 580226 285368 584960 285424
rect 580165 285366 584960 285368
rect 580165 285363 580231 285366
rect 583520 285276 584960 285366
rect 580165 284474 580231 284477
rect 576350 284472 580231 284474
rect 576350 284416 580170 284472
rect 580226 284416 580231 284472
rect 576350 284414 580231 284416
rect 576350 284398 576410 284414
rect 580165 284411 580231 284414
rect 575920 284338 576410 284398
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 3417 279030 3483 279033
rect 3417 279028 4048 279030
rect 3417 278972 3422 279028
rect 3478 278972 4048 279028
rect 3417 278970 4048 278972
rect 3417 278967 3483 278970
rect 579613 272234 579679 272237
rect 583520 272234 584960 272324
rect 579613 272232 584960 272234
rect 579613 272176 579618 272232
rect 579674 272176 584960 272232
rect 579613 272174 584960 272176
rect 579613 272171 579679 272174
rect 583520 272084 584960 272174
rect 579521 271146 579587 271149
rect 576350 271144 579587 271146
rect 576350 271100 579526 271144
rect 575920 271088 579526 271100
rect 579582 271088 579587 271144
rect 575920 271086 579587 271088
rect 575920 271040 576410 271086
rect 579521 271083 579587 271086
rect -960 267202 480 267292
rect 3417 267202 3483 267205
rect -960 267200 3483 267202
rect -960 267144 3422 267200
rect 3478 267144 3483 267200
rect -960 267142 3483 267144
rect -960 267052 480 267142
rect 3417 267139 3483 267142
rect 3417 265976 3483 265979
rect 3417 265974 4048 265976
rect 3417 265918 3422 265974
rect 3478 265918 4048 265974
rect 3417 265916 4048 265918
rect 3417 265913 3483 265916
rect 580901 258906 580967 258909
rect 583520 258906 584960 258996
rect 580901 258904 584960 258906
rect 580901 258848 580906 258904
rect 580962 258848 584960 258904
rect 580901 258846 584960 258848
rect 580901 258843 580967 258846
rect 583520 258756 584960 258846
rect 578877 257682 578943 257685
rect 576350 257680 578943 257682
rect 575920 257624 578882 257680
rect 578938 257624 578943 257680
rect 575920 257622 578943 257624
rect 575920 257620 576410 257622
rect 578877 257619 578943 257622
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 3417 252800 3483 252803
rect 3417 252798 4048 252800
rect 3417 252742 3422 252798
rect 3478 252742 4048 252798
rect 3417 252740 4048 252742
rect 3417 252737 3483 252740
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 580165 244490 580231 244493
rect 576350 244488 580231 244490
rect 576350 244432 580170 244488
rect 580226 244432 580231 244488
rect 576350 244430 580231 244432
rect 576350 244382 576410 244430
rect 580165 244427 580231 244430
rect 575920 244322 576410 244382
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 3417 239746 3483 239749
rect 3417 239744 4048 239746
rect 3417 239688 3422 239744
rect 3478 239688 4048 239744
rect 3417 239686 4048 239688
rect 3417 239683 3483 239686
rect 579613 232386 579679 232389
rect 583520 232386 584960 232476
rect 579613 232384 584960 232386
rect 579613 232328 579618 232384
rect 579674 232328 584960 232384
rect 579613 232326 584960 232328
rect 579613 232323 579679 232326
rect 583520 232236 584960 232326
rect 579521 231162 579587 231165
rect 576350 231160 579587 231162
rect 576350 231104 579526 231160
rect 579582 231104 579587 231160
rect 576350 231102 579587 231104
rect 576350 231084 576410 231102
rect 579521 231099 579587 231102
rect 575920 231024 576410 231084
rect -960 228034 480 228124
rect 3417 228034 3483 228037
rect -960 228032 3483 228034
rect -960 227976 3422 228032
rect 3478 227976 3483 228032
rect -960 227974 3483 227976
rect -960 227884 480 227974
rect 3417 227971 3483 227974
rect 3417 226692 3483 226695
rect 3417 226690 4048 226692
rect 3417 226634 3422 226690
rect 3478 226634 4048 226690
rect 3417 226632 4048 226634
rect 3417 226629 3483 226632
rect 579613 219058 579679 219061
rect 583520 219058 584960 219148
rect 579613 219056 584960 219058
rect 579613 219000 579618 219056
rect 579674 219000 584960 219056
rect 579613 218998 584960 219000
rect 579613 218995 579679 218998
rect 583520 218908 584960 218998
rect 579521 217698 579587 217701
rect 576350 217696 579587 217698
rect 576350 217664 579526 217696
rect 575920 217640 579526 217664
rect 579582 217640 579587 217696
rect 575920 217638 579587 217640
rect 575920 217604 576410 217638
rect 579521 217635 579587 217638
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 3417 213516 3483 213519
rect 3417 213514 4048 213516
rect 3417 213458 3422 213514
rect 3478 213458 4048 213514
rect 3417 213456 4048 213458
rect 3417 213453 3483 213456
rect 579613 205730 579679 205733
rect 583520 205730 584960 205820
rect 579613 205728 584960 205730
rect 579613 205672 579618 205728
rect 579674 205672 584960 205728
rect 579613 205670 584960 205672
rect 579613 205667 579679 205670
rect 583520 205580 584960 205670
rect 579521 204370 579587 204373
rect 576350 204368 579587 204370
rect 576350 204366 579526 204368
rect 575920 204312 579526 204366
rect 579582 204312 579587 204368
rect 575920 204310 579587 204312
rect 575920 204306 576410 204310
rect 579521 204307 579587 204310
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 3417 200462 3483 200465
rect 3417 200460 4048 200462
rect 3417 200404 3422 200460
rect 3478 200404 4048 200460
rect 3417 200402 4048 200404
rect 3417 200399 3483 200402
rect 579613 192538 579679 192541
rect 583520 192538 584960 192628
rect 579613 192536 584960 192538
rect 579613 192480 579618 192536
rect 579674 192480 584960 192536
rect 579613 192478 584960 192480
rect 579613 192475 579679 192478
rect 583520 192388 584960 192478
rect 575920 191042 576410 191068
rect 579521 191042 579587 191045
rect 575920 191040 579587 191042
rect 575920 191008 579526 191040
rect 576350 190984 579526 191008
rect 579582 190984 579587 191040
rect 576350 190982 579587 190984
rect 579521 190979 579587 190982
rect -960 188866 480 188956
rect 3601 188866 3667 188869
rect -960 188864 3667 188866
rect -960 188808 3606 188864
rect 3662 188808 3667 188864
rect -960 188806 3667 188808
rect -960 188716 480 188806
rect 3601 188803 3667 188806
rect 3601 187408 3667 187411
rect 3601 187406 4048 187408
rect 3601 187350 3606 187406
rect 3662 187350 4048 187406
rect 3601 187348 4048 187350
rect 3601 187345 3667 187348
rect 579613 179210 579679 179213
rect 583520 179210 584960 179300
rect 579613 179208 584960 179210
rect 579613 179152 579618 179208
rect 579674 179152 584960 179208
rect 579613 179150 584960 179152
rect 579613 179147 579679 179150
rect 583520 179060 584960 179150
rect 579521 177714 579587 177717
rect 576350 177712 579587 177714
rect 576350 177656 579526 177712
rect 579582 177656 579587 177712
rect 576350 177654 579587 177656
rect 576350 177648 576410 177654
rect 579521 177651 579587 177654
rect 575920 177588 576410 177648
rect -960 175946 480 176036
rect 3417 175946 3483 175949
rect -960 175944 3483 175946
rect -960 175888 3422 175944
rect 3478 175888 3483 175944
rect -960 175886 3483 175888
rect -960 175796 480 175886
rect 3417 175883 3483 175886
rect 3417 174232 3483 174235
rect 3417 174230 4048 174232
rect 3417 174174 3422 174230
rect 3478 174174 4048 174230
rect 3417 174172 4048 174174
rect 3417 174169 3483 174172
rect 579613 165882 579679 165885
rect 583520 165882 584960 165972
rect 579613 165880 584960 165882
rect 579613 165824 579618 165880
rect 579674 165824 584960 165880
rect 579613 165822 584960 165824
rect 579613 165819 579679 165822
rect 583520 165732 584960 165822
rect 579521 164386 579587 164389
rect 576350 164384 579587 164386
rect 576350 164350 579526 164384
rect 575920 164328 579526 164350
rect 579582 164328 579587 164384
rect 575920 164326 579587 164328
rect 575920 164290 576410 164326
rect 579521 164323 579587 164326
rect -960 162890 480 162980
rect 2129 162890 2195 162893
rect -960 162888 2195 162890
rect -960 162832 2134 162888
rect 2190 162832 2195 162888
rect -960 162830 2195 162832
rect -960 162740 480 162830
rect 2129 162827 2195 162830
rect 2129 161122 2195 161125
rect 3374 161122 4048 161178
rect 2129 161120 4048 161122
rect 2129 161064 2134 161120
rect 2190 161118 4048 161120
rect 2190 161064 3434 161118
rect 2129 161062 3434 161064
rect 2129 161059 2195 161062
rect 580901 152690 580967 152693
rect 583520 152690 584960 152780
rect 580901 152688 584960 152690
rect 580901 152632 580906 152688
rect 580962 152632 584960 152688
rect 580901 152630 584960 152632
rect 580901 152627 580967 152630
rect 583520 152540 584960 152630
rect 578509 151058 578575 151061
rect 576350 151056 578575 151058
rect 576350 151052 578514 151056
rect 575920 151000 578514 151052
rect 578570 151000 578575 151056
rect 575920 150998 578575 151000
rect 575920 150992 576410 150998
rect 578509 150995 578575 150998
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 3417 148124 3483 148127
rect 3417 148122 4048 148124
rect 3417 148066 3422 148122
rect 3478 148066 4048 148122
rect 3417 148064 4048 148066
rect 3417 148061 3483 148064
rect 579613 139362 579679 139365
rect 583520 139362 584960 139452
rect 579613 139360 584960 139362
rect 579613 139304 579618 139360
rect 579674 139304 584960 139360
rect 579613 139302 584960 139304
rect 579613 139299 579679 139302
rect 583520 139212 584960 139302
rect 575920 137594 576410 137632
rect 579521 137594 579587 137597
rect 575920 137592 579587 137594
rect 575920 137572 579526 137592
rect 576350 137536 579526 137572
rect 579582 137536 579587 137592
rect 576350 137534 579587 137536
rect 579521 137531 579587 137534
rect -960 136778 480 136868
rect 2129 136778 2195 136781
rect -960 136776 2195 136778
rect -960 136720 2134 136776
rect 2190 136720 2195 136776
rect -960 136718 2195 136720
rect -960 136628 480 136718
rect 2129 136715 2195 136718
rect 2129 135010 2195 135013
rect 3374 135010 4048 135070
rect 2129 135008 3434 135010
rect 2129 134952 2134 135008
rect 2190 134952 3434 135008
rect 2129 134950 3434 134952
rect 2129 134947 2195 134950
rect 579613 126034 579679 126037
rect 583520 126034 584960 126124
rect 579613 126032 584960 126034
rect 579613 125976 579618 126032
rect 579674 125976 584960 126032
rect 579613 125974 584960 125976
rect 579613 125971 579679 125974
rect 583520 125884 584960 125974
rect 579521 124402 579587 124405
rect 576350 124400 579587 124402
rect 576350 124344 579526 124400
rect 579582 124344 579587 124400
rect 576350 124342 579587 124344
rect 576350 124334 576410 124342
rect 579521 124339 579587 124342
rect 575920 124274 576410 124334
rect -960 123722 480 123812
rect 3417 123722 3483 123725
rect -960 123720 3483 123722
rect -960 123664 3422 123720
rect 3478 123664 3483 123720
rect -960 123662 3483 123664
rect -960 123572 480 123662
rect 3417 123659 3483 123662
rect 3417 121894 3483 121897
rect 3417 121892 4048 121894
rect 3417 121836 3422 121892
rect 3478 121836 4048 121892
rect 3417 121834 4048 121836
rect 3417 121831 3483 121834
rect 579613 112842 579679 112845
rect 583520 112842 584960 112932
rect 579613 112840 584960 112842
rect 579613 112784 579618 112840
rect 579674 112784 584960 112840
rect 579613 112782 584960 112784
rect 579613 112779 579679 112782
rect 583520 112692 584960 112782
rect 579521 110938 579587 110941
rect 576350 110936 579587 110938
rect 576350 110914 579526 110936
rect 575920 110880 579526 110914
rect 579582 110880 579587 110936
rect 575920 110878 579587 110880
rect 575920 110854 576410 110878
rect 579521 110875 579587 110878
rect -960 110666 480 110756
rect 2129 110666 2195 110669
rect -960 110664 2195 110666
rect -960 110608 2134 110664
rect 2190 110608 2195 110664
rect -960 110606 2195 110608
rect -960 110516 480 110606
rect 2129 110603 2195 110606
rect 2129 108898 2195 108901
rect 2129 108896 3434 108898
rect 2129 108840 2134 108896
rect 2190 108840 3434 108896
rect 2129 108838 4048 108840
rect 2129 108835 2195 108838
rect 3374 108780 4048 108838
rect 579613 99514 579679 99517
rect 583520 99514 584960 99604
rect 579613 99512 584960 99514
rect 579613 99456 579618 99512
rect 579674 99456 584960 99512
rect 579613 99454 584960 99456
rect 579613 99451 579679 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect 575920 97610 576410 97616
rect 579521 97610 579587 97613
rect 575920 97608 579587 97610
rect 575920 97556 579526 97608
rect -960 97550 3483 97552
rect 576350 97552 579526 97556
rect 579582 97552 579587 97608
rect 576350 97550 579587 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 579521 97547 579587 97550
rect 3417 95786 3483 95789
rect 3417 95784 4048 95786
rect 3417 95728 3422 95784
rect 3478 95728 4048 95784
rect 3417 95726 4048 95728
rect 3417 95723 3483 95726
rect 579613 86186 579679 86189
rect 583520 86186 584960 86276
rect 579613 86184 584960 86186
rect 579613 86128 579618 86184
rect 579674 86128 584960 86184
rect 579613 86126 584960 86128
rect 579613 86123 579679 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 2129 84690 2195 84693
rect -960 84688 2195 84690
rect -960 84632 2134 84688
rect 2190 84632 2195 84688
rect -960 84630 2195 84632
rect -960 84540 480 84630
rect 2129 84627 2195 84630
rect 575920 84282 576410 84318
rect 579521 84282 579587 84285
rect 575920 84280 579587 84282
rect 575920 84258 579526 84280
rect 576350 84224 579526 84258
rect 579582 84224 579587 84280
rect 576350 84222 579587 84224
rect 579521 84219 579587 84222
rect 2129 82650 2195 82653
rect 2129 82648 3434 82650
rect 2129 82592 2134 82648
rect 2190 82610 3434 82648
rect 2190 82592 4048 82610
rect 2129 82590 4048 82592
rect 2129 82587 2195 82590
rect 3374 82550 4048 82590
rect 579613 72994 579679 72997
rect 583520 72994 584960 73084
rect 579613 72992 584960 72994
rect 579613 72936 579618 72992
rect 579674 72936 584960 72992
rect 579613 72934 584960 72936
rect 579613 72931 579679 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 579521 70954 579587 70957
rect 576350 70952 579587 70954
rect 576350 70898 579526 70952
rect 575920 70896 579526 70898
rect 579582 70896 579587 70952
rect 575920 70894 579587 70896
rect 575920 70838 576410 70894
rect 579521 70891 579587 70894
rect 3417 69556 3483 69559
rect 3417 69554 4048 69556
rect 3417 69498 3422 69554
rect 3478 69498 4048 69554
rect 3417 69496 4048 69498
rect 3417 69493 3483 69496
rect 579613 59666 579679 59669
rect 583520 59666 584960 59756
rect 579613 59664 584960 59666
rect 579613 59608 579618 59664
rect 579674 59608 584960 59664
rect 579613 59606 584960 59608
rect 579613 59603 579679 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2129 58578 2195 58581
rect -960 58576 2195 58578
rect -960 58520 2134 58576
rect 2190 58520 2195 58576
rect -960 58518 2195 58520
rect -960 58428 480 58518
rect 2129 58515 2195 58518
rect 579521 57626 579587 57629
rect 576350 57624 579587 57626
rect 576350 57600 579526 57624
rect 575920 57568 579526 57600
rect 579582 57568 579587 57624
rect 575920 57566 579587 57568
rect 575920 57540 576410 57566
rect 579521 57563 579587 57566
rect 2129 56538 2195 56541
rect 2129 56536 3434 56538
rect 2129 56480 2134 56536
rect 2190 56502 3434 56536
rect 2190 56480 4048 56502
rect 2129 56478 4048 56480
rect 2129 56475 2195 56478
rect 3374 56442 4048 56478
rect 579981 46338 580047 46341
rect 583520 46338 584960 46428
rect 579981 46336 584960 46338
rect 579981 46280 579986 46336
rect 580042 46280 584960 46336
rect 579981 46278 584960 46280
rect 579981 46275 580047 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 575920 44298 576410 44302
rect 578325 44298 578391 44301
rect 575920 44296 578391 44298
rect 575920 44242 578330 44296
rect 576350 44240 578330 44242
rect 578386 44240 578391 44296
rect 576350 44238 578391 44240
rect 578325 44235 578391 44238
rect 3417 43326 3483 43329
rect 3417 43324 4048 43326
rect 3417 43268 3422 43324
rect 3478 43268 4048 43324
rect 3417 43266 4048 43268
rect 3417 43263 3483 43266
rect 579613 33146 579679 33149
rect 583520 33146 584960 33236
rect 579613 33144 584960 33146
rect 579613 33088 579618 33144
rect 579674 33088 584960 33144
rect 579613 33086 584960 33088
rect 579613 33083 579679 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2129 32466 2195 32469
rect -960 32464 2195 32466
rect -960 32408 2134 32464
rect 2190 32408 2195 32464
rect -960 32406 2195 32408
rect -960 32316 480 32406
rect 2129 32403 2195 32406
rect 579521 30970 579587 30973
rect 576350 30968 579587 30970
rect 576350 30912 579526 30968
rect 579582 30912 579587 30968
rect 576350 30910 579587 30912
rect 576350 30882 576410 30910
rect 579521 30907 579587 30910
rect 575920 30822 576410 30882
rect 2129 30290 2195 30293
rect 2129 30288 3434 30290
rect 2129 30232 2134 30288
rect 2190 30272 3434 30288
rect 2190 30232 4048 30272
rect 2129 30230 4048 30232
rect 2129 30227 2195 30230
rect 3374 30212 4048 30230
rect 579613 19818 579679 19821
rect 583520 19818 584960 19908
rect 579613 19816 584960 19818
rect 579613 19760 579618 19816
rect 579674 19760 584960 19816
rect 579613 19758 584960 19760
rect 579613 19755 579679 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 2037 19410 2103 19413
rect -960 19408 2103 19410
rect -960 19352 2042 19408
rect 2098 19352 2103 19408
rect -960 19350 2103 19352
rect -960 19260 480 19350
rect 2037 19347 2103 19350
rect 579521 17642 579587 17645
rect 576350 17640 579587 17642
rect 576350 17584 579526 17640
rect 579582 17584 579587 17640
rect 575920 17582 579587 17584
rect 575920 17524 576410 17582
rect 579521 17579 579587 17582
rect 2037 17234 2103 17237
rect 2037 17232 3434 17234
rect 2037 17176 2042 17232
rect 2098 17218 3434 17232
rect 2098 17176 4048 17218
rect 2037 17174 4048 17176
rect 2037 17171 2103 17174
rect 3374 17158 4048 17174
rect 579613 6626 579679 6629
rect 583520 6626 584960 6716
rect 579613 6624 584960 6626
rect -960 6490 480 6580
rect 579613 6568 579618 6624
rect 579674 6568 584960 6624
rect 579613 6566 584960 6568
rect 579613 6563 579679 6566
rect 2773 6490 2839 6493
rect -960 6488 2839 6490
rect -960 6432 2778 6488
rect 2834 6432 2839 6488
rect 583520 6476 584960 6566
rect -960 6430 2839 6432
rect -960 6340 480 6430
rect 2773 6427 2839 6430
rect 2773 4178 2839 4181
rect 579521 4178 579587 4181
rect 2773 4176 3802 4178
rect 2773 4120 2778 4176
rect 2834 4164 3802 4176
rect 576166 4176 579587 4178
rect 576166 4164 579526 4176
rect 2834 4120 4048 4164
rect 2773 4118 4048 4120
rect 2773 4115 2839 4118
rect 3742 4104 4048 4118
rect 575920 4120 579526 4164
rect 579582 4120 579587 4176
rect 575920 4118 579587 4120
rect 575920 4104 576226 4118
rect 579521 4115 579587 4118
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 700008 2414 704282
rect 5514 700008 6134 706202
rect 9234 700008 9854 708122
rect 12954 700008 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 700008 20414 705242
rect 23514 700008 24134 707162
rect 27234 700008 27854 709082
rect 30954 700008 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 700008 38414 704282
rect 41514 700008 42134 706202
rect 45234 700008 45854 708122
rect 48954 700008 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 700008 56414 705242
rect 59514 700008 60134 707162
rect 63234 700008 63854 709082
rect 66954 700008 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 700008 74414 704282
rect 77514 700008 78134 706202
rect 81234 700008 81854 708122
rect 84954 700008 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 700008 92414 705242
rect 95514 700008 96134 707162
rect 99234 700008 99854 709082
rect 102954 700008 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 700008 110414 704282
rect 113514 700008 114134 706202
rect 117234 700008 117854 708122
rect 120954 700008 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 700008 128414 705242
rect 131514 700008 132134 707162
rect 135234 700008 135854 709082
rect 138954 700008 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 700008 146414 704282
rect 149514 700008 150134 706202
rect 153234 700008 153854 708122
rect 156954 700008 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 700008 164414 705242
rect 167514 700008 168134 707162
rect 171234 700008 171854 709082
rect 174954 700008 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 700008 182414 704282
rect 185514 700008 186134 706202
rect 189234 700008 189854 708122
rect 192954 700008 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 700008 200414 705242
rect 203514 700008 204134 707162
rect 207234 700008 207854 709082
rect 210954 700008 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 700008 218414 704282
rect 221514 700008 222134 706202
rect 225234 700008 225854 708122
rect 228954 700008 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 700008 236414 705242
rect 239514 700008 240134 707162
rect 243234 700008 243854 709082
rect 246954 700008 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 700008 254414 704282
rect 257514 700008 258134 706202
rect 261234 700008 261854 708122
rect 264954 700008 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 700008 272414 705242
rect 275514 700008 276134 707162
rect 279234 700008 279854 709082
rect 282954 700008 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 700008 290414 704282
rect 293514 700008 294134 706202
rect 297234 700008 297854 708122
rect 300954 700008 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 700008 308414 705242
rect 311514 700008 312134 707162
rect 315234 700008 315854 709082
rect 318954 700008 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 700008 326414 704282
rect 329514 700008 330134 706202
rect 333234 700008 333854 708122
rect 336954 700008 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 700008 344414 705242
rect 347514 700008 348134 707162
rect 351234 700008 351854 709082
rect 354954 700008 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 700008 362414 704282
rect 365514 700008 366134 706202
rect 369234 700008 369854 708122
rect 372954 700008 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 700008 380414 705242
rect 383514 700008 384134 707162
rect 387234 700008 387854 709082
rect 390954 700008 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 700008 398414 704282
rect 401514 700008 402134 706202
rect 405234 700008 405854 708122
rect 408954 700008 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 700008 416414 705242
rect 419514 700008 420134 707162
rect 423234 700008 423854 709082
rect 426954 700008 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 700008 434414 704282
rect 437514 700008 438134 706202
rect 441234 700008 441854 708122
rect 444954 700008 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 700008 452414 705242
rect 455514 700008 456134 707162
rect 459234 700008 459854 709082
rect 462954 700008 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 700008 470414 704282
rect 473514 700008 474134 706202
rect 477234 700008 477854 708122
rect 480954 700008 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 700008 488414 705242
rect 491514 700008 492134 707162
rect 495234 700008 495854 709082
rect 498954 700008 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 700008 506414 704282
rect 509514 700008 510134 706202
rect 513234 700008 513854 708122
rect 516954 700008 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 700008 524414 705242
rect 527514 700008 528134 707162
rect 531234 700008 531854 709082
rect 534954 700008 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 700008 542414 704282
rect 545514 700008 546134 706202
rect 549234 700008 549854 708122
rect 552954 700008 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 700008 560414 705242
rect 563514 700008 564134 707162
rect 567234 700008 567854 709082
rect 570954 700008 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 700008 578414 704282
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect 9084 687454 9704 687486
rect 9084 687218 9116 687454
rect 9352 687218 9436 687454
rect 9672 687218 9704 687454
rect 9084 687134 9704 687218
rect 9084 686898 9116 687134
rect 9352 686898 9436 687134
rect 9672 686898 9704 687134
rect 9084 686866 9704 686898
rect 56620 687454 57240 687486
rect 56620 687218 56652 687454
rect 56888 687218 56972 687454
rect 57208 687218 57240 687454
rect 56620 687134 57240 687218
rect 56620 686898 56652 687134
rect 56888 686898 56972 687134
rect 57208 686898 57240 687134
rect 56620 686866 57240 686898
rect 92620 687454 93240 687486
rect 92620 687218 92652 687454
rect 92888 687218 92972 687454
rect 93208 687218 93240 687454
rect 92620 687134 93240 687218
rect 92620 686898 92652 687134
rect 92888 686898 92972 687134
rect 93208 686898 93240 687134
rect 92620 686866 93240 686898
rect 128620 687454 129240 687486
rect 128620 687218 128652 687454
rect 128888 687218 128972 687454
rect 129208 687218 129240 687454
rect 128620 687134 129240 687218
rect 128620 686898 128652 687134
rect 128888 686898 128972 687134
rect 129208 686898 129240 687134
rect 128620 686866 129240 686898
rect 164620 687454 165240 687486
rect 164620 687218 164652 687454
rect 164888 687218 164972 687454
rect 165208 687218 165240 687454
rect 164620 687134 165240 687218
rect 164620 686898 164652 687134
rect 164888 686898 164972 687134
rect 165208 686898 165240 687134
rect 164620 686866 165240 686898
rect 200620 687454 201240 687486
rect 200620 687218 200652 687454
rect 200888 687218 200972 687454
rect 201208 687218 201240 687454
rect 200620 687134 201240 687218
rect 200620 686898 200652 687134
rect 200888 686898 200972 687134
rect 201208 686898 201240 687134
rect 200620 686866 201240 686898
rect 236620 687454 237240 687486
rect 236620 687218 236652 687454
rect 236888 687218 236972 687454
rect 237208 687218 237240 687454
rect 236620 687134 237240 687218
rect 236620 686898 236652 687134
rect 236888 686898 236972 687134
rect 237208 686898 237240 687134
rect 236620 686866 237240 686898
rect 272620 687454 273240 687486
rect 272620 687218 272652 687454
rect 272888 687218 272972 687454
rect 273208 687218 273240 687454
rect 272620 687134 273240 687218
rect 272620 686898 272652 687134
rect 272888 686898 272972 687134
rect 273208 686898 273240 687134
rect 272620 686866 273240 686898
rect 308620 687454 309240 687486
rect 308620 687218 308652 687454
rect 308888 687218 308972 687454
rect 309208 687218 309240 687454
rect 308620 687134 309240 687218
rect 308620 686898 308652 687134
rect 308888 686898 308972 687134
rect 309208 686898 309240 687134
rect 308620 686866 309240 686898
rect 344620 687454 345240 687486
rect 344620 687218 344652 687454
rect 344888 687218 344972 687454
rect 345208 687218 345240 687454
rect 344620 687134 345240 687218
rect 344620 686898 344652 687134
rect 344888 686898 344972 687134
rect 345208 686898 345240 687134
rect 344620 686866 345240 686898
rect 380620 687454 381240 687486
rect 380620 687218 380652 687454
rect 380888 687218 380972 687454
rect 381208 687218 381240 687454
rect 380620 687134 381240 687218
rect 380620 686898 380652 687134
rect 380888 686898 380972 687134
rect 381208 686898 381240 687134
rect 380620 686866 381240 686898
rect 416620 687454 417240 687486
rect 416620 687218 416652 687454
rect 416888 687218 416972 687454
rect 417208 687218 417240 687454
rect 416620 687134 417240 687218
rect 416620 686898 416652 687134
rect 416888 686898 416972 687134
rect 417208 686898 417240 687134
rect 416620 686866 417240 686898
rect 452620 687454 453240 687486
rect 452620 687218 452652 687454
rect 452888 687218 452972 687454
rect 453208 687218 453240 687454
rect 452620 687134 453240 687218
rect 452620 686898 452652 687134
rect 452888 686898 452972 687134
rect 453208 686898 453240 687134
rect 452620 686866 453240 686898
rect 488620 687454 489240 687486
rect 488620 687218 488652 687454
rect 488888 687218 488972 687454
rect 489208 687218 489240 687454
rect 488620 687134 489240 687218
rect 488620 686898 488652 687134
rect 488888 686898 488972 687134
rect 489208 686898 489240 687134
rect 488620 686866 489240 686898
rect 524620 687454 525240 687486
rect 524620 687218 524652 687454
rect 524888 687218 524972 687454
rect 525208 687218 525240 687454
rect 524620 687134 525240 687218
rect 524620 686898 524652 687134
rect 524888 686898 524972 687134
rect 525208 686898 525240 687134
rect 524620 686866 525240 686898
rect 560620 687454 561240 687486
rect 560620 687218 560652 687454
rect 560888 687218 560972 687454
rect 561208 687218 561240 687454
rect 560620 687134 561240 687218
rect 560620 686898 560652 687134
rect 560888 686898 560972 687134
rect 561208 686898 561240 687134
rect 560620 686866 561240 686898
rect 570260 687454 570880 687486
rect 570260 687218 570292 687454
rect 570528 687218 570612 687454
rect 570848 687218 570880 687454
rect 570260 687134 570880 687218
rect 570260 686898 570292 687134
rect 570528 686898 570612 687134
rect 570848 686898 570880 687134
rect 570260 686866 570880 686898
rect 7844 669454 8464 669486
rect 7844 669218 7876 669454
rect 8112 669218 8196 669454
rect 8432 669218 8464 669454
rect 7844 669134 8464 669218
rect 7844 668898 7876 669134
rect 8112 668898 8196 669134
rect 8432 668898 8464 669134
rect 7844 668866 8464 668898
rect 38000 669454 38620 669486
rect 38000 669218 38032 669454
rect 38268 669218 38352 669454
rect 38588 669218 38620 669454
rect 38000 669134 38620 669218
rect 38000 668898 38032 669134
rect 38268 668898 38352 669134
rect 38588 668898 38620 669134
rect 38000 668866 38620 668898
rect 74000 669454 74620 669486
rect 74000 669218 74032 669454
rect 74268 669218 74352 669454
rect 74588 669218 74620 669454
rect 74000 669134 74620 669218
rect 74000 668898 74032 669134
rect 74268 668898 74352 669134
rect 74588 668898 74620 669134
rect 74000 668866 74620 668898
rect 100381 669454 100741 669486
rect 100381 669218 100443 669454
rect 100679 669218 100741 669454
rect 100381 669134 100741 669218
rect 100381 668898 100443 669134
rect 100679 668898 100741 669134
rect 100381 668866 100741 668898
rect 198857 669454 199217 669486
rect 198857 669218 198919 669454
rect 199155 669218 199217 669454
rect 198857 669134 199217 669218
rect 198857 668898 198919 669134
rect 199155 668898 199217 669134
rect 198857 668866 199217 668898
rect 216337 669454 216697 669486
rect 216337 669218 216399 669454
rect 216635 669218 216697 669454
rect 216337 669134 216697 669218
rect 216337 668898 216399 669134
rect 216635 668898 216697 669134
rect 216337 668866 216697 668898
rect 314813 669454 315173 669486
rect 314813 669218 314875 669454
rect 315111 669218 315173 669454
rect 314813 669134 315173 669218
rect 314813 668898 314875 669134
rect 315111 668898 315173 669134
rect 314813 668866 315173 668898
rect 326000 669454 326620 669486
rect 326000 669218 326032 669454
rect 326268 669218 326352 669454
rect 326588 669218 326620 669454
rect 326000 669134 326620 669218
rect 326000 668898 326032 669134
rect 326268 668898 326352 669134
rect 326588 668898 326620 669134
rect 326000 668866 326620 668898
rect 332293 669454 332653 669486
rect 332293 669218 332355 669454
rect 332591 669218 332653 669454
rect 332293 669134 332653 669218
rect 332293 668898 332355 669134
rect 332591 668898 332653 669134
rect 332293 668866 332653 668898
rect 430769 669454 431129 669486
rect 430769 669218 430831 669454
rect 431067 669218 431129 669454
rect 430769 669134 431129 669218
rect 430769 668898 430831 669134
rect 431067 668898 431129 669134
rect 430769 668866 431129 668898
rect 434000 669454 434620 669486
rect 434000 669218 434032 669454
rect 434268 669218 434352 669454
rect 434588 669218 434620 669454
rect 434000 669134 434620 669218
rect 434000 668898 434032 669134
rect 434268 668898 434352 669134
rect 434588 668898 434620 669134
rect 434000 668866 434620 668898
rect 448249 669454 448609 669486
rect 448249 669218 448311 669454
rect 448547 669218 448609 669454
rect 448249 669134 448609 669218
rect 448249 668898 448311 669134
rect 448547 668898 448609 669134
rect 448249 668866 448609 668898
rect 546725 669454 547085 669486
rect 546725 669218 546787 669454
rect 547023 669218 547085 669454
rect 546725 669134 547085 669218
rect 546725 668898 546787 669134
rect 547023 668898 547085 669134
rect 546725 668866 547085 668898
rect 571500 669454 572120 669486
rect 571500 669218 571532 669454
rect 571768 669218 571852 669454
rect 572088 669218 572120 669454
rect 571500 669134 572120 669218
rect 571500 668898 571532 669134
rect 571768 668898 571852 669134
rect 572088 668898 572120 669134
rect 571500 668866 572120 668898
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect 9084 651454 9704 651486
rect 9084 651218 9116 651454
rect 9352 651218 9436 651454
rect 9672 651218 9704 651454
rect 9084 651134 9704 651218
rect 9084 650898 9116 651134
rect 9352 650898 9436 651134
rect 9672 650898 9704 651134
rect 9084 650866 9704 650898
rect 56620 651454 57240 651486
rect 56620 651218 56652 651454
rect 56888 651218 56972 651454
rect 57208 651218 57240 651454
rect 56620 651134 57240 651218
rect 56620 650898 56652 651134
rect 56888 650898 56972 651134
rect 57208 650898 57240 651134
rect 56620 650866 57240 650898
rect 92620 651454 93240 651486
rect 92620 651218 92652 651454
rect 92888 651218 92972 651454
rect 93208 651218 93240 651454
rect 92620 651134 93240 651218
rect 92620 650898 92652 651134
rect 92888 650898 92972 651134
rect 93208 650898 93240 651134
rect 92620 650866 93240 650898
rect 101101 651454 101461 651486
rect 101101 651218 101163 651454
rect 101399 651218 101461 651454
rect 101101 651134 101461 651218
rect 101101 650898 101163 651134
rect 101399 650898 101461 651134
rect 101101 650866 101461 650898
rect 198137 651454 198497 651486
rect 198137 651218 198199 651454
rect 198435 651218 198497 651454
rect 198137 651134 198497 651218
rect 198137 650898 198199 651134
rect 198435 650898 198497 651134
rect 198137 650866 198497 650898
rect 200620 651454 201240 651486
rect 200620 651218 200652 651454
rect 200888 651218 200972 651454
rect 201208 651218 201240 651454
rect 200620 651134 201240 651218
rect 200620 650898 200652 651134
rect 200888 650898 200972 651134
rect 201208 650898 201240 651134
rect 200620 650866 201240 650898
rect 217057 651454 217417 651486
rect 217057 651218 217119 651454
rect 217355 651218 217417 651454
rect 217057 651134 217417 651218
rect 217057 650898 217119 651134
rect 217355 650898 217417 651134
rect 217057 650866 217417 650898
rect 314093 651454 314453 651486
rect 314093 651218 314155 651454
rect 314391 651218 314453 651454
rect 314093 651134 314453 651218
rect 314093 650898 314155 651134
rect 314391 650898 314453 651134
rect 314093 650866 314453 650898
rect 333013 651454 333373 651486
rect 333013 651218 333075 651454
rect 333311 651218 333373 651454
rect 333013 651134 333373 651218
rect 333013 650898 333075 651134
rect 333311 650898 333373 651134
rect 333013 650866 333373 650898
rect 430049 651454 430409 651486
rect 430049 651218 430111 651454
rect 430347 651218 430409 651454
rect 430049 651134 430409 651218
rect 430049 650898 430111 651134
rect 430347 650898 430409 651134
rect 430049 650866 430409 650898
rect 448969 651454 449329 651486
rect 448969 651218 449031 651454
rect 449267 651218 449329 651454
rect 448969 651134 449329 651218
rect 448969 650898 449031 651134
rect 449267 650898 449329 651134
rect 448969 650866 449329 650898
rect 546005 651454 546365 651486
rect 546005 651218 546067 651454
rect 546303 651218 546365 651454
rect 546005 651134 546365 651218
rect 546005 650898 546067 651134
rect 546303 650898 546365 651134
rect 546005 650866 546365 650898
rect 560620 651454 561240 651486
rect 560620 651218 560652 651454
rect 560888 651218 560972 651454
rect 561208 651218 561240 651454
rect 560620 651134 561240 651218
rect 560620 650898 560652 651134
rect 560888 650898 560972 651134
rect 561208 650898 561240 651134
rect 560620 650866 561240 650898
rect 570260 651454 570880 651486
rect 570260 651218 570292 651454
rect 570528 651218 570612 651454
rect 570848 651218 570880 651454
rect 570260 651134 570880 651218
rect 570260 650898 570292 651134
rect 570528 650898 570612 651134
rect 570848 650898 570880 651134
rect 570260 650866 570880 650898
rect 7844 633454 8464 633486
rect 7844 633218 7876 633454
rect 8112 633218 8196 633454
rect 8432 633218 8464 633454
rect 7844 633134 8464 633218
rect 7844 632898 7876 633134
rect 8112 632898 8196 633134
rect 8432 632898 8464 633134
rect 7844 632866 8464 632898
rect 38000 633454 38620 633486
rect 38000 633218 38032 633454
rect 38268 633218 38352 633454
rect 38588 633218 38620 633454
rect 38000 633134 38620 633218
rect 38000 632898 38032 633134
rect 38268 632898 38352 633134
rect 38588 632898 38620 633134
rect 38000 632866 38620 632898
rect 74000 633454 74620 633486
rect 74000 633218 74032 633454
rect 74268 633218 74352 633454
rect 74588 633218 74620 633454
rect 74000 633134 74620 633218
rect 74000 632898 74032 633134
rect 74268 632898 74352 633134
rect 74588 632898 74620 633134
rect 74000 632866 74620 632898
rect 100381 633454 100741 633486
rect 100381 633218 100443 633454
rect 100679 633218 100741 633454
rect 100381 633134 100741 633218
rect 100381 632898 100443 633134
rect 100679 632898 100741 633134
rect 100381 632866 100741 632898
rect 198857 633454 199217 633486
rect 198857 633218 198919 633454
rect 199155 633218 199217 633454
rect 198857 633134 199217 633218
rect 198857 632898 198919 633134
rect 199155 632898 199217 633134
rect 198857 632866 199217 632898
rect 216337 633454 216697 633486
rect 216337 633218 216399 633454
rect 216635 633218 216697 633454
rect 216337 633134 216697 633218
rect 216337 632898 216399 633134
rect 216635 632898 216697 633134
rect 216337 632866 216697 632898
rect 314813 633454 315173 633486
rect 314813 633218 314875 633454
rect 315111 633218 315173 633454
rect 314813 633134 315173 633218
rect 314813 632898 314875 633134
rect 315111 632898 315173 633134
rect 314813 632866 315173 632898
rect 326000 633454 326620 633486
rect 326000 633218 326032 633454
rect 326268 633218 326352 633454
rect 326588 633218 326620 633454
rect 326000 633134 326620 633218
rect 326000 632898 326032 633134
rect 326268 632898 326352 633134
rect 326588 632898 326620 633134
rect 326000 632866 326620 632898
rect 332293 633454 332653 633486
rect 332293 633218 332355 633454
rect 332591 633218 332653 633454
rect 332293 633134 332653 633218
rect 332293 632898 332355 633134
rect 332591 632898 332653 633134
rect 332293 632866 332653 632898
rect 430769 633454 431129 633486
rect 430769 633218 430831 633454
rect 431067 633218 431129 633454
rect 430769 633134 431129 633218
rect 430769 632898 430831 633134
rect 431067 632898 431129 633134
rect 430769 632866 431129 632898
rect 434000 633454 434620 633486
rect 434000 633218 434032 633454
rect 434268 633218 434352 633454
rect 434588 633218 434620 633454
rect 434000 633134 434620 633218
rect 434000 632898 434032 633134
rect 434268 632898 434352 633134
rect 434588 632898 434620 633134
rect 434000 632866 434620 632898
rect 448249 633454 448609 633486
rect 448249 633218 448311 633454
rect 448547 633218 448609 633454
rect 448249 633134 448609 633218
rect 448249 632898 448311 633134
rect 448547 632898 448609 633134
rect 448249 632866 448609 632898
rect 546725 633454 547085 633486
rect 546725 633218 546787 633454
rect 547023 633218 547085 633454
rect 546725 633134 547085 633218
rect 546725 632898 546787 633134
rect 547023 632898 547085 633134
rect 546725 632866 547085 632898
rect 571500 633454 572120 633486
rect 571500 633218 571532 633454
rect 571768 633218 571852 633454
rect 572088 633218 572120 633454
rect 571500 633134 572120 633218
rect 571500 632898 571532 633134
rect 571768 632898 571852 633134
rect 572088 632898 572120 633134
rect 571500 632866 572120 632898
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect 9084 615454 9704 615486
rect 9084 615218 9116 615454
rect 9352 615218 9436 615454
rect 9672 615218 9704 615454
rect 9084 615134 9704 615218
rect 9084 614898 9116 615134
rect 9352 614898 9436 615134
rect 9672 614898 9704 615134
rect 9084 614866 9704 614898
rect 56620 615454 57240 615486
rect 56620 615218 56652 615454
rect 56888 615218 56972 615454
rect 57208 615218 57240 615454
rect 56620 615134 57240 615218
rect 56620 614898 56652 615134
rect 56888 614898 56972 615134
rect 57208 614898 57240 615134
rect 56620 614866 57240 614898
rect 92620 615454 93240 615486
rect 92620 615218 92652 615454
rect 92888 615218 92972 615454
rect 93208 615218 93240 615454
rect 92620 615134 93240 615218
rect 92620 614898 92652 615134
rect 92888 614898 92972 615134
rect 93208 614898 93240 615134
rect 92620 614866 93240 614898
rect 101101 615454 101461 615486
rect 101101 615218 101163 615454
rect 101399 615218 101461 615454
rect 101101 615134 101461 615218
rect 101101 614898 101163 615134
rect 101399 614898 101461 615134
rect 101101 614866 101461 614898
rect 198137 615454 198497 615486
rect 198137 615218 198199 615454
rect 198435 615218 198497 615454
rect 198137 615134 198497 615218
rect 198137 614898 198199 615134
rect 198435 614898 198497 615134
rect 198137 614866 198497 614898
rect 200620 615454 201240 615486
rect 200620 615218 200652 615454
rect 200888 615218 200972 615454
rect 201208 615218 201240 615454
rect 200620 615134 201240 615218
rect 200620 614898 200652 615134
rect 200888 614898 200972 615134
rect 201208 614898 201240 615134
rect 200620 614866 201240 614898
rect 217057 615454 217417 615486
rect 217057 615218 217119 615454
rect 217355 615218 217417 615454
rect 217057 615134 217417 615218
rect 217057 614898 217119 615134
rect 217355 614898 217417 615134
rect 217057 614866 217417 614898
rect 314093 615454 314453 615486
rect 314093 615218 314155 615454
rect 314391 615218 314453 615454
rect 314093 615134 314453 615218
rect 314093 614898 314155 615134
rect 314391 614898 314453 615134
rect 314093 614866 314453 614898
rect 333013 615454 333373 615486
rect 333013 615218 333075 615454
rect 333311 615218 333373 615454
rect 333013 615134 333373 615218
rect 333013 614898 333075 615134
rect 333311 614898 333373 615134
rect 333013 614866 333373 614898
rect 430049 615454 430409 615486
rect 430049 615218 430111 615454
rect 430347 615218 430409 615454
rect 430049 615134 430409 615218
rect 430049 614898 430111 615134
rect 430347 614898 430409 615134
rect 430049 614866 430409 614898
rect 448969 615454 449329 615486
rect 448969 615218 449031 615454
rect 449267 615218 449329 615454
rect 448969 615134 449329 615218
rect 448969 614898 449031 615134
rect 449267 614898 449329 615134
rect 448969 614866 449329 614898
rect 546005 615454 546365 615486
rect 546005 615218 546067 615454
rect 546303 615218 546365 615454
rect 546005 615134 546365 615218
rect 546005 614898 546067 615134
rect 546303 614898 546365 615134
rect 546005 614866 546365 614898
rect 560620 615454 561240 615486
rect 560620 615218 560652 615454
rect 560888 615218 560972 615454
rect 561208 615218 561240 615454
rect 560620 615134 561240 615218
rect 560620 614898 560652 615134
rect 560888 614898 560972 615134
rect 561208 614898 561240 615134
rect 560620 614866 561240 614898
rect 570260 615454 570880 615486
rect 570260 615218 570292 615454
rect 570528 615218 570612 615454
rect 570848 615218 570880 615454
rect 570260 615134 570880 615218
rect 570260 614898 570292 615134
rect 570528 614898 570612 615134
rect 570848 614898 570880 615134
rect 570260 614866 570880 614898
rect 7844 597454 8464 597486
rect 7844 597218 7876 597454
rect 8112 597218 8196 597454
rect 8432 597218 8464 597454
rect 7844 597134 8464 597218
rect 7844 596898 7876 597134
rect 8112 596898 8196 597134
rect 8432 596898 8464 597134
rect 7844 596866 8464 596898
rect 38000 597454 38620 597486
rect 38000 597218 38032 597454
rect 38268 597218 38352 597454
rect 38588 597218 38620 597454
rect 38000 597134 38620 597218
rect 38000 596898 38032 597134
rect 38268 596898 38352 597134
rect 38588 596898 38620 597134
rect 38000 596866 38620 596898
rect 74000 597454 74620 597486
rect 74000 597218 74032 597454
rect 74268 597218 74352 597454
rect 74588 597218 74620 597454
rect 74000 597134 74620 597218
rect 74000 596898 74032 597134
rect 74268 596898 74352 597134
rect 74588 596898 74620 597134
rect 74000 596866 74620 596898
rect 100381 597454 100741 597486
rect 100381 597218 100443 597454
rect 100679 597218 100741 597454
rect 100381 597134 100741 597218
rect 100381 596898 100443 597134
rect 100679 596898 100741 597134
rect 100381 596866 100741 596898
rect 198857 597454 199217 597486
rect 198857 597218 198919 597454
rect 199155 597218 199217 597454
rect 198857 597134 199217 597218
rect 198857 596898 198919 597134
rect 199155 596898 199217 597134
rect 198857 596866 199217 596898
rect 216337 597454 216697 597486
rect 216337 597218 216399 597454
rect 216635 597218 216697 597454
rect 216337 597134 216697 597218
rect 216337 596898 216399 597134
rect 216635 596898 216697 597134
rect 216337 596866 216697 596898
rect 314813 597454 315173 597486
rect 314813 597218 314875 597454
rect 315111 597218 315173 597454
rect 314813 597134 315173 597218
rect 314813 596898 314875 597134
rect 315111 596898 315173 597134
rect 314813 596866 315173 596898
rect 326000 597454 326620 597486
rect 326000 597218 326032 597454
rect 326268 597218 326352 597454
rect 326588 597218 326620 597454
rect 326000 597134 326620 597218
rect 326000 596898 326032 597134
rect 326268 596898 326352 597134
rect 326588 596898 326620 597134
rect 326000 596866 326620 596898
rect 332293 597454 332653 597486
rect 332293 597218 332355 597454
rect 332591 597218 332653 597454
rect 332293 597134 332653 597218
rect 332293 596898 332355 597134
rect 332591 596898 332653 597134
rect 332293 596866 332653 596898
rect 430769 597454 431129 597486
rect 430769 597218 430831 597454
rect 431067 597218 431129 597454
rect 430769 597134 431129 597218
rect 430769 596898 430831 597134
rect 431067 596898 431129 597134
rect 430769 596866 431129 596898
rect 434000 597454 434620 597486
rect 434000 597218 434032 597454
rect 434268 597218 434352 597454
rect 434588 597218 434620 597454
rect 434000 597134 434620 597218
rect 434000 596898 434032 597134
rect 434268 596898 434352 597134
rect 434588 596898 434620 597134
rect 434000 596866 434620 596898
rect 448249 597454 448609 597486
rect 448249 597218 448311 597454
rect 448547 597218 448609 597454
rect 448249 597134 448609 597218
rect 448249 596898 448311 597134
rect 448547 596898 448609 597134
rect 448249 596866 448609 596898
rect 546725 597454 547085 597486
rect 546725 597218 546787 597454
rect 547023 597218 547085 597454
rect 546725 597134 547085 597218
rect 546725 596898 546787 597134
rect 547023 596898 547085 597134
rect 546725 596866 547085 596898
rect 571500 597454 572120 597486
rect 571500 597218 571532 597454
rect 571768 597218 571852 597454
rect 572088 597218 572120 597454
rect 571500 597134 572120 597218
rect 571500 596898 571532 597134
rect 571768 596898 571852 597134
rect 572088 596898 572120 597134
rect 571500 596866 572120 596898
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect 9084 579454 9704 579486
rect 9084 579218 9116 579454
rect 9352 579218 9436 579454
rect 9672 579218 9704 579454
rect 9084 579134 9704 579218
rect 9084 578898 9116 579134
rect 9352 578898 9436 579134
rect 9672 578898 9704 579134
rect 9084 578866 9704 578898
rect 56620 579454 57240 579486
rect 56620 579218 56652 579454
rect 56888 579218 56972 579454
rect 57208 579218 57240 579454
rect 56620 579134 57240 579218
rect 56620 578898 56652 579134
rect 56888 578898 56972 579134
rect 57208 578898 57240 579134
rect 56620 578866 57240 578898
rect 92620 579454 93240 579486
rect 92620 579218 92652 579454
rect 92888 579218 92972 579454
rect 93208 579218 93240 579454
rect 92620 579134 93240 579218
rect 92620 578898 92652 579134
rect 92888 578898 92972 579134
rect 93208 578898 93240 579134
rect 92620 578866 93240 578898
rect 128620 579454 129240 579486
rect 128620 579218 128652 579454
rect 128888 579218 128972 579454
rect 129208 579218 129240 579454
rect 128620 579134 129240 579218
rect 128620 578898 128652 579134
rect 128888 578898 128972 579134
rect 129208 578898 129240 579134
rect 128620 578866 129240 578898
rect 164620 579454 165240 579486
rect 164620 579218 164652 579454
rect 164888 579218 164972 579454
rect 165208 579218 165240 579454
rect 164620 579134 165240 579218
rect 164620 578898 164652 579134
rect 164888 578898 164972 579134
rect 165208 578898 165240 579134
rect 164620 578866 165240 578898
rect 200620 579454 201240 579486
rect 200620 579218 200652 579454
rect 200888 579218 200972 579454
rect 201208 579218 201240 579454
rect 200620 579134 201240 579218
rect 200620 578898 200652 579134
rect 200888 578898 200972 579134
rect 201208 578898 201240 579134
rect 200620 578866 201240 578898
rect 236620 579454 237240 579486
rect 236620 579218 236652 579454
rect 236888 579218 236972 579454
rect 237208 579218 237240 579454
rect 236620 579134 237240 579218
rect 236620 578898 236652 579134
rect 236888 578898 236972 579134
rect 237208 578898 237240 579134
rect 236620 578866 237240 578898
rect 272620 579454 273240 579486
rect 272620 579218 272652 579454
rect 272888 579218 272972 579454
rect 273208 579218 273240 579454
rect 272620 579134 273240 579218
rect 272620 578898 272652 579134
rect 272888 578898 272972 579134
rect 273208 578898 273240 579134
rect 272620 578866 273240 578898
rect 308620 579454 309240 579486
rect 308620 579218 308652 579454
rect 308888 579218 308972 579454
rect 309208 579218 309240 579454
rect 308620 579134 309240 579218
rect 308620 578898 308652 579134
rect 308888 578898 308972 579134
rect 309208 578898 309240 579134
rect 308620 578866 309240 578898
rect 344620 579454 345240 579486
rect 344620 579218 344652 579454
rect 344888 579218 344972 579454
rect 345208 579218 345240 579454
rect 344620 579134 345240 579218
rect 344620 578898 344652 579134
rect 344888 578898 344972 579134
rect 345208 578898 345240 579134
rect 344620 578866 345240 578898
rect 380620 579454 381240 579486
rect 380620 579218 380652 579454
rect 380888 579218 380972 579454
rect 381208 579218 381240 579454
rect 380620 579134 381240 579218
rect 380620 578898 380652 579134
rect 380888 578898 380972 579134
rect 381208 578898 381240 579134
rect 380620 578866 381240 578898
rect 416620 579454 417240 579486
rect 416620 579218 416652 579454
rect 416888 579218 416972 579454
rect 417208 579218 417240 579454
rect 416620 579134 417240 579218
rect 416620 578898 416652 579134
rect 416888 578898 416972 579134
rect 417208 578898 417240 579134
rect 416620 578866 417240 578898
rect 452620 579454 453240 579486
rect 452620 579218 452652 579454
rect 452888 579218 452972 579454
rect 453208 579218 453240 579454
rect 452620 579134 453240 579218
rect 452620 578898 452652 579134
rect 452888 578898 452972 579134
rect 453208 578898 453240 579134
rect 452620 578866 453240 578898
rect 488620 579454 489240 579486
rect 488620 579218 488652 579454
rect 488888 579218 488972 579454
rect 489208 579218 489240 579454
rect 488620 579134 489240 579218
rect 488620 578898 488652 579134
rect 488888 578898 488972 579134
rect 489208 578898 489240 579134
rect 488620 578866 489240 578898
rect 524620 579454 525240 579486
rect 524620 579218 524652 579454
rect 524888 579218 524972 579454
rect 525208 579218 525240 579454
rect 524620 579134 525240 579218
rect 524620 578898 524652 579134
rect 524888 578898 524972 579134
rect 525208 578898 525240 579134
rect 524620 578866 525240 578898
rect 560620 579454 561240 579486
rect 560620 579218 560652 579454
rect 560888 579218 560972 579454
rect 561208 579218 561240 579454
rect 560620 579134 561240 579218
rect 560620 578898 560652 579134
rect 560888 578898 560972 579134
rect 561208 578898 561240 579134
rect 560620 578866 561240 578898
rect 570260 579454 570880 579486
rect 570260 579218 570292 579454
rect 570528 579218 570612 579454
rect 570848 579218 570880 579454
rect 570260 579134 570880 579218
rect 570260 578898 570292 579134
rect 570528 578898 570612 579134
rect 570848 578898 570880 579134
rect 570260 578866 570880 578898
rect 7844 561454 8464 561486
rect 7844 561218 7876 561454
rect 8112 561218 8196 561454
rect 8432 561218 8464 561454
rect 7844 561134 8464 561218
rect 7844 560898 7876 561134
rect 8112 560898 8196 561134
rect 8432 560898 8464 561134
rect 7844 560866 8464 560898
rect 38000 561454 38620 561486
rect 38000 561218 38032 561454
rect 38268 561218 38352 561454
rect 38588 561218 38620 561454
rect 38000 561134 38620 561218
rect 38000 560898 38032 561134
rect 38268 560898 38352 561134
rect 38588 560898 38620 561134
rect 38000 560866 38620 560898
rect 74000 561454 74620 561486
rect 74000 561218 74032 561454
rect 74268 561218 74352 561454
rect 74588 561218 74620 561454
rect 74000 561134 74620 561218
rect 74000 560898 74032 561134
rect 74268 560898 74352 561134
rect 74588 560898 74620 561134
rect 74000 560866 74620 560898
rect 110000 561454 110620 561486
rect 110000 561218 110032 561454
rect 110268 561218 110352 561454
rect 110588 561218 110620 561454
rect 110000 561134 110620 561218
rect 110000 560898 110032 561134
rect 110268 560898 110352 561134
rect 110588 560898 110620 561134
rect 110000 560866 110620 560898
rect 146000 561454 146620 561486
rect 146000 561218 146032 561454
rect 146268 561218 146352 561454
rect 146588 561218 146620 561454
rect 146000 561134 146620 561218
rect 146000 560898 146032 561134
rect 146268 560898 146352 561134
rect 146588 560898 146620 561134
rect 146000 560866 146620 560898
rect 182000 561454 182620 561486
rect 182000 561218 182032 561454
rect 182268 561218 182352 561454
rect 182588 561218 182620 561454
rect 182000 561134 182620 561218
rect 182000 560898 182032 561134
rect 182268 560898 182352 561134
rect 182588 560898 182620 561134
rect 182000 560866 182620 560898
rect 218000 561454 218620 561486
rect 218000 561218 218032 561454
rect 218268 561218 218352 561454
rect 218588 561218 218620 561454
rect 218000 561134 218620 561218
rect 218000 560898 218032 561134
rect 218268 560898 218352 561134
rect 218588 560898 218620 561134
rect 218000 560866 218620 560898
rect 254000 561454 254620 561486
rect 254000 561218 254032 561454
rect 254268 561218 254352 561454
rect 254588 561218 254620 561454
rect 254000 561134 254620 561218
rect 254000 560898 254032 561134
rect 254268 560898 254352 561134
rect 254588 560898 254620 561134
rect 254000 560866 254620 560898
rect 290000 561454 290620 561486
rect 290000 561218 290032 561454
rect 290268 561218 290352 561454
rect 290588 561218 290620 561454
rect 290000 561134 290620 561218
rect 290000 560898 290032 561134
rect 290268 560898 290352 561134
rect 290588 560898 290620 561134
rect 290000 560866 290620 560898
rect 326000 561454 326620 561486
rect 326000 561218 326032 561454
rect 326268 561218 326352 561454
rect 326588 561218 326620 561454
rect 326000 561134 326620 561218
rect 326000 560898 326032 561134
rect 326268 560898 326352 561134
rect 326588 560898 326620 561134
rect 326000 560866 326620 560898
rect 332293 561454 332653 561486
rect 332293 561218 332355 561454
rect 332591 561218 332653 561454
rect 332293 561134 332653 561218
rect 332293 560898 332355 561134
rect 332591 560898 332653 561134
rect 332293 560866 332653 560898
rect 430769 561454 431129 561486
rect 430769 561218 430831 561454
rect 431067 561218 431129 561454
rect 430769 561134 431129 561218
rect 430769 560898 430831 561134
rect 431067 560898 431129 561134
rect 430769 560866 431129 560898
rect 434000 561454 434620 561486
rect 434000 561218 434032 561454
rect 434268 561218 434352 561454
rect 434588 561218 434620 561454
rect 434000 561134 434620 561218
rect 434000 560898 434032 561134
rect 434268 560898 434352 561134
rect 434588 560898 434620 561134
rect 434000 560866 434620 560898
rect 448249 561454 448609 561486
rect 448249 561218 448311 561454
rect 448547 561218 448609 561454
rect 448249 561134 448609 561218
rect 448249 560898 448311 561134
rect 448547 560898 448609 561134
rect 448249 560866 448609 560898
rect 546725 561454 547085 561486
rect 546725 561218 546787 561454
rect 547023 561218 547085 561454
rect 546725 561134 547085 561218
rect 546725 560898 546787 561134
rect 547023 560898 547085 561134
rect 546725 560866 547085 560898
rect 571500 561454 572120 561486
rect 571500 561218 571532 561454
rect 571768 561218 571852 561454
rect 572088 561218 572120 561454
rect 571500 561134 572120 561218
rect 571500 560898 571532 561134
rect 571768 560898 571852 561134
rect 572088 560898 572120 561134
rect 571500 560866 572120 560898
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect 9084 543454 9704 543486
rect 9084 543218 9116 543454
rect 9352 543218 9436 543454
rect 9672 543218 9704 543454
rect 9084 543134 9704 543218
rect 9084 542898 9116 543134
rect 9352 542898 9436 543134
rect 9672 542898 9704 543134
rect 9084 542866 9704 542898
rect 56620 543454 57240 543486
rect 56620 543218 56652 543454
rect 56888 543218 56972 543454
rect 57208 543218 57240 543454
rect 56620 543134 57240 543218
rect 56620 542898 56652 543134
rect 56888 542898 56972 543134
rect 57208 542898 57240 543134
rect 56620 542866 57240 542898
rect 92620 543454 93240 543486
rect 92620 543218 92652 543454
rect 92888 543218 92972 543454
rect 93208 543218 93240 543454
rect 92620 543134 93240 543218
rect 92620 542898 92652 543134
rect 92888 542898 92972 543134
rect 93208 542898 93240 543134
rect 92620 542866 93240 542898
rect 128620 543454 129240 543486
rect 128620 543218 128652 543454
rect 128888 543218 128972 543454
rect 129208 543218 129240 543454
rect 128620 543134 129240 543218
rect 128620 542898 128652 543134
rect 128888 542898 128972 543134
rect 129208 542898 129240 543134
rect 128620 542866 129240 542898
rect 164620 543454 165240 543486
rect 164620 543218 164652 543454
rect 164888 543218 164972 543454
rect 165208 543218 165240 543454
rect 164620 543134 165240 543218
rect 164620 542898 164652 543134
rect 164888 542898 164972 543134
rect 165208 542898 165240 543134
rect 164620 542866 165240 542898
rect 200620 543454 201240 543486
rect 200620 543218 200652 543454
rect 200888 543218 200972 543454
rect 201208 543218 201240 543454
rect 200620 543134 201240 543218
rect 200620 542898 200652 543134
rect 200888 542898 200972 543134
rect 201208 542898 201240 543134
rect 200620 542866 201240 542898
rect 236620 543454 237240 543486
rect 236620 543218 236652 543454
rect 236888 543218 236972 543454
rect 237208 543218 237240 543454
rect 236620 543134 237240 543218
rect 236620 542898 236652 543134
rect 236888 542898 236972 543134
rect 237208 542898 237240 543134
rect 236620 542866 237240 542898
rect 272620 543454 273240 543486
rect 272620 543218 272652 543454
rect 272888 543218 272972 543454
rect 273208 543218 273240 543454
rect 272620 543134 273240 543218
rect 272620 542898 272652 543134
rect 272888 542898 272972 543134
rect 273208 542898 273240 543134
rect 272620 542866 273240 542898
rect 308620 543454 309240 543486
rect 308620 543218 308652 543454
rect 308888 543218 308972 543454
rect 309208 543218 309240 543454
rect 308620 543134 309240 543218
rect 308620 542898 308652 543134
rect 308888 542898 308972 543134
rect 309208 542898 309240 543134
rect 308620 542866 309240 542898
rect 333013 543454 333373 543486
rect 333013 543218 333075 543454
rect 333311 543218 333373 543454
rect 333013 543134 333373 543218
rect 333013 542898 333075 543134
rect 333311 542898 333373 543134
rect 333013 542866 333373 542898
rect 430049 543454 430409 543486
rect 430049 543218 430111 543454
rect 430347 543218 430409 543454
rect 430049 543134 430409 543218
rect 430049 542898 430111 543134
rect 430347 542898 430409 543134
rect 430049 542866 430409 542898
rect 448969 543454 449329 543486
rect 448969 543218 449031 543454
rect 449267 543218 449329 543454
rect 448969 543134 449329 543218
rect 448969 542898 449031 543134
rect 449267 542898 449329 543134
rect 448969 542866 449329 542898
rect 546005 543454 546365 543486
rect 546005 543218 546067 543454
rect 546303 543218 546365 543454
rect 546005 543134 546365 543218
rect 546005 542898 546067 543134
rect 546303 542898 546365 543134
rect 546005 542866 546365 542898
rect 560620 543454 561240 543486
rect 560620 543218 560652 543454
rect 560888 543218 560972 543454
rect 561208 543218 561240 543454
rect 560620 543134 561240 543218
rect 560620 542898 560652 543134
rect 560888 542898 560972 543134
rect 561208 542898 561240 543134
rect 560620 542866 561240 542898
rect 570260 543454 570880 543486
rect 570260 543218 570292 543454
rect 570528 543218 570612 543454
rect 570848 543218 570880 543454
rect 570260 543134 570880 543218
rect 570260 542898 570292 543134
rect 570528 542898 570612 543134
rect 570848 542898 570880 543134
rect 570260 542866 570880 542898
rect 7844 525454 8464 525486
rect 7844 525218 7876 525454
rect 8112 525218 8196 525454
rect 8432 525218 8464 525454
rect 7844 525134 8464 525218
rect 7844 524898 7876 525134
rect 8112 524898 8196 525134
rect 8432 524898 8464 525134
rect 7844 524866 8464 524898
rect 38000 525454 38620 525486
rect 38000 525218 38032 525454
rect 38268 525218 38352 525454
rect 38588 525218 38620 525454
rect 38000 525134 38620 525218
rect 38000 524898 38032 525134
rect 38268 524898 38352 525134
rect 38588 524898 38620 525134
rect 38000 524866 38620 524898
rect 74000 525454 74620 525486
rect 74000 525218 74032 525454
rect 74268 525218 74352 525454
rect 74588 525218 74620 525454
rect 74000 525134 74620 525218
rect 74000 524898 74032 525134
rect 74268 524898 74352 525134
rect 74588 524898 74620 525134
rect 74000 524866 74620 524898
rect 110000 525454 110620 525486
rect 110000 525218 110032 525454
rect 110268 525218 110352 525454
rect 110588 525218 110620 525454
rect 110000 525134 110620 525218
rect 110000 524898 110032 525134
rect 110268 524898 110352 525134
rect 110588 524898 110620 525134
rect 110000 524866 110620 524898
rect 146000 525454 146620 525486
rect 146000 525218 146032 525454
rect 146268 525218 146352 525454
rect 146588 525218 146620 525454
rect 146000 525134 146620 525218
rect 146000 524898 146032 525134
rect 146268 524898 146352 525134
rect 146588 524898 146620 525134
rect 146000 524866 146620 524898
rect 182000 525454 182620 525486
rect 182000 525218 182032 525454
rect 182268 525218 182352 525454
rect 182588 525218 182620 525454
rect 182000 525134 182620 525218
rect 182000 524898 182032 525134
rect 182268 524898 182352 525134
rect 182588 524898 182620 525134
rect 182000 524866 182620 524898
rect 218000 525454 218620 525486
rect 218000 525218 218032 525454
rect 218268 525218 218352 525454
rect 218588 525218 218620 525454
rect 218000 525134 218620 525218
rect 218000 524898 218032 525134
rect 218268 524898 218352 525134
rect 218588 524898 218620 525134
rect 218000 524866 218620 524898
rect 254000 525454 254620 525486
rect 254000 525218 254032 525454
rect 254268 525218 254352 525454
rect 254588 525218 254620 525454
rect 254000 525134 254620 525218
rect 254000 524898 254032 525134
rect 254268 524898 254352 525134
rect 254588 524898 254620 525134
rect 254000 524866 254620 524898
rect 290000 525454 290620 525486
rect 290000 525218 290032 525454
rect 290268 525218 290352 525454
rect 290588 525218 290620 525454
rect 290000 525134 290620 525218
rect 290000 524898 290032 525134
rect 290268 524898 290352 525134
rect 290588 524898 290620 525134
rect 290000 524866 290620 524898
rect 326000 525454 326620 525486
rect 326000 525218 326032 525454
rect 326268 525218 326352 525454
rect 326588 525218 326620 525454
rect 326000 525134 326620 525218
rect 326000 524898 326032 525134
rect 326268 524898 326352 525134
rect 326588 524898 326620 525134
rect 326000 524866 326620 524898
rect 332293 525454 332653 525486
rect 332293 525218 332355 525454
rect 332591 525218 332653 525454
rect 332293 525134 332653 525218
rect 332293 524898 332355 525134
rect 332591 524898 332653 525134
rect 332293 524866 332653 524898
rect 430769 525454 431129 525486
rect 430769 525218 430831 525454
rect 431067 525218 431129 525454
rect 430769 525134 431129 525218
rect 430769 524898 430831 525134
rect 431067 524898 431129 525134
rect 430769 524866 431129 524898
rect 434000 525454 434620 525486
rect 434000 525218 434032 525454
rect 434268 525218 434352 525454
rect 434588 525218 434620 525454
rect 434000 525134 434620 525218
rect 434000 524898 434032 525134
rect 434268 524898 434352 525134
rect 434588 524898 434620 525134
rect 434000 524866 434620 524898
rect 448249 525454 448609 525486
rect 448249 525218 448311 525454
rect 448547 525218 448609 525454
rect 448249 525134 448609 525218
rect 448249 524898 448311 525134
rect 448547 524898 448609 525134
rect 448249 524866 448609 524898
rect 546725 525454 547085 525486
rect 546725 525218 546787 525454
rect 547023 525218 547085 525454
rect 546725 525134 547085 525218
rect 546725 524898 546787 525134
rect 547023 524898 547085 525134
rect 546725 524866 547085 524898
rect 571500 525454 572120 525486
rect 571500 525218 571532 525454
rect 571768 525218 571852 525454
rect 572088 525218 572120 525454
rect 571500 525134 572120 525218
rect 571500 524898 571532 525134
rect 571768 524898 571852 525134
rect 572088 524898 572120 525134
rect 571500 524866 572120 524898
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect 9084 507454 9704 507486
rect 9084 507218 9116 507454
rect 9352 507218 9436 507454
rect 9672 507218 9704 507454
rect 9084 507134 9704 507218
rect 9084 506898 9116 507134
rect 9352 506898 9436 507134
rect 9672 506898 9704 507134
rect 9084 506866 9704 506898
rect 56620 507454 57240 507486
rect 56620 507218 56652 507454
rect 56888 507218 56972 507454
rect 57208 507218 57240 507454
rect 56620 507134 57240 507218
rect 56620 506898 56652 507134
rect 56888 506898 56972 507134
rect 57208 506898 57240 507134
rect 56620 506866 57240 506898
rect 92620 507454 93240 507486
rect 92620 507218 92652 507454
rect 92888 507218 92972 507454
rect 93208 507218 93240 507454
rect 92620 507134 93240 507218
rect 92620 506898 92652 507134
rect 92888 506898 92972 507134
rect 93208 506898 93240 507134
rect 92620 506866 93240 506898
rect 128620 507454 129240 507486
rect 128620 507218 128652 507454
rect 128888 507218 128972 507454
rect 129208 507218 129240 507454
rect 128620 507134 129240 507218
rect 128620 506898 128652 507134
rect 128888 506898 128972 507134
rect 129208 506898 129240 507134
rect 128620 506866 129240 506898
rect 164620 507454 165240 507486
rect 164620 507218 164652 507454
rect 164888 507218 164972 507454
rect 165208 507218 165240 507454
rect 164620 507134 165240 507218
rect 164620 506898 164652 507134
rect 164888 506898 164972 507134
rect 165208 506898 165240 507134
rect 164620 506866 165240 506898
rect 200620 507454 201240 507486
rect 200620 507218 200652 507454
rect 200888 507218 200972 507454
rect 201208 507218 201240 507454
rect 200620 507134 201240 507218
rect 200620 506898 200652 507134
rect 200888 506898 200972 507134
rect 201208 506898 201240 507134
rect 200620 506866 201240 506898
rect 236620 507454 237240 507486
rect 236620 507218 236652 507454
rect 236888 507218 236972 507454
rect 237208 507218 237240 507454
rect 236620 507134 237240 507218
rect 236620 506898 236652 507134
rect 236888 506898 236972 507134
rect 237208 506898 237240 507134
rect 236620 506866 237240 506898
rect 272620 507454 273240 507486
rect 272620 507218 272652 507454
rect 272888 507218 272972 507454
rect 273208 507218 273240 507454
rect 272620 507134 273240 507218
rect 272620 506898 272652 507134
rect 272888 506898 272972 507134
rect 273208 506898 273240 507134
rect 272620 506866 273240 506898
rect 308620 507454 309240 507486
rect 308620 507218 308652 507454
rect 308888 507218 308972 507454
rect 309208 507218 309240 507454
rect 308620 507134 309240 507218
rect 308620 506898 308652 507134
rect 308888 506898 308972 507134
rect 309208 506898 309240 507134
rect 308620 506866 309240 506898
rect 333013 507454 333373 507486
rect 333013 507218 333075 507454
rect 333311 507218 333373 507454
rect 333013 507134 333373 507218
rect 333013 506898 333075 507134
rect 333311 506898 333373 507134
rect 333013 506866 333373 506898
rect 430049 507454 430409 507486
rect 430049 507218 430111 507454
rect 430347 507218 430409 507454
rect 430049 507134 430409 507218
rect 430049 506898 430111 507134
rect 430347 506898 430409 507134
rect 430049 506866 430409 506898
rect 448969 507454 449329 507486
rect 448969 507218 449031 507454
rect 449267 507218 449329 507454
rect 448969 507134 449329 507218
rect 448969 506898 449031 507134
rect 449267 506898 449329 507134
rect 448969 506866 449329 506898
rect 546005 507454 546365 507486
rect 546005 507218 546067 507454
rect 546303 507218 546365 507454
rect 546005 507134 546365 507218
rect 546005 506898 546067 507134
rect 546303 506898 546365 507134
rect 546005 506866 546365 506898
rect 560620 507454 561240 507486
rect 560620 507218 560652 507454
rect 560888 507218 560972 507454
rect 561208 507218 561240 507454
rect 560620 507134 561240 507218
rect 560620 506898 560652 507134
rect 560888 506898 560972 507134
rect 561208 506898 561240 507134
rect 560620 506866 561240 506898
rect 570260 507454 570880 507486
rect 570260 507218 570292 507454
rect 570528 507218 570612 507454
rect 570848 507218 570880 507454
rect 570260 507134 570880 507218
rect 570260 506898 570292 507134
rect 570528 506898 570612 507134
rect 570848 506898 570880 507134
rect 570260 506866 570880 506898
rect 7844 489454 8464 489486
rect 7844 489218 7876 489454
rect 8112 489218 8196 489454
rect 8432 489218 8464 489454
rect 7844 489134 8464 489218
rect 7844 488898 7876 489134
rect 8112 488898 8196 489134
rect 8432 488898 8464 489134
rect 7844 488866 8464 488898
rect 38000 489454 38620 489486
rect 38000 489218 38032 489454
rect 38268 489218 38352 489454
rect 38588 489218 38620 489454
rect 38000 489134 38620 489218
rect 38000 488898 38032 489134
rect 38268 488898 38352 489134
rect 38588 488898 38620 489134
rect 38000 488866 38620 488898
rect 74000 489454 74620 489486
rect 74000 489218 74032 489454
rect 74268 489218 74352 489454
rect 74588 489218 74620 489454
rect 74000 489134 74620 489218
rect 74000 488898 74032 489134
rect 74268 488898 74352 489134
rect 74588 488898 74620 489134
rect 74000 488866 74620 488898
rect 110000 489454 110620 489486
rect 110000 489218 110032 489454
rect 110268 489218 110352 489454
rect 110588 489218 110620 489454
rect 110000 489134 110620 489218
rect 110000 488898 110032 489134
rect 110268 488898 110352 489134
rect 110588 488898 110620 489134
rect 110000 488866 110620 488898
rect 146000 489454 146620 489486
rect 146000 489218 146032 489454
rect 146268 489218 146352 489454
rect 146588 489218 146620 489454
rect 146000 489134 146620 489218
rect 146000 488898 146032 489134
rect 146268 488898 146352 489134
rect 146588 488898 146620 489134
rect 146000 488866 146620 488898
rect 182000 489454 182620 489486
rect 182000 489218 182032 489454
rect 182268 489218 182352 489454
rect 182588 489218 182620 489454
rect 182000 489134 182620 489218
rect 182000 488898 182032 489134
rect 182268 488898 182352 489134
rect 182588 488898 182620 489134
rect 182000 488866 182620 488898
rect 218000 489454 218620 489486
rect 218000 489218 218032 489454
rect 218268 489218 218352 489454
rect 218588 489218 218620 489454
rect 218000 489134 218620 489218
rect 218000 488898 218032 489134
rect 218268 488898 218352 489134
rect 218588 488898 218620 489134
rect 218000 488866 218620 488898
rect 254000 489454 254620 489486
rect 254000 489218 254032 489454
rect 254268 489218 254352 489454
rect 254588 489218 254620 489454
rect 254000 489134 254620 489218
rect 254000 488898 254032 489134
rect 254268 488898 254352 489134
rect 254588 488898 254620 489134
rect 254000 488866 254620 488898
rect 290000 489454 290620 489486
rect 290000 489218 290032 489454
rect 290268 489218 290352 489454
rect 290588 489218 290620 489454
rect 290000 489134 290620 489218
rect 290000 488898 290032 489134
rect 290268 488898 290352 489134
rect 290588 488898 290620 489134
rect 290000 488866 290620 488898
rect 326000 489454 326620 489486
rect 326000 489218 326032 489454
rect 326268 489218 326352 489454
rect 326588 489218 326620 489454
rect 326000 489134 326620 489218
rect 326000 488898 326032 489134
rect 326268 488898 326352 489134
rect 326588 488898 326620 489134
rect 326000 488866 326620 488898
rect 362000 489454 362620 489486
rect 362000 489218 362032 489454
rect 362268 489218 362352 489454
rect 362588 489218 362620 489454
rect 362000 489134 362620 489218
rect 362000 488898 362032 489134
rect 362268 488898 362352 489134
rect 362588 488898 362620 489134
rect 362000 488866 362620 488898
rect 398000 489454 398620 489486
rect 398000 489218 398032 489454
rect 398268 489218 398352 489454
rect 398588 489218 398620 489454
rect 398000 489134 398620 489218
rect 398000 488898 398032 489134
rect 398268 488898 398352 489134
rect 398588 488898 398620 489134
rect 398000 488866 398620 488898
rect 434000 489454 434620 489486
rect 434000 489218 434032 489454
rect 434268 489218 434352 489454
rect 434588 489218 434620 489454
rect 434000 489134 434620 489218
rect 434000 488898 434032 489134
rect 434268 488898 434352 489134
rect 434588 488898 434620 489134
rect 434000 488866 434620 488898
rect 470000 489454 470620 489486
rect 470000 489218 470032 489454
rect 470268 489218 470352 489454
rect 470588 489218 470620 489454
rect 470000 489134 470620 489218
rect 470000 488898 470032 489134
rect 470268 488898 470352 489134
rect 470588 488898 470620 489134
rect 470000 488866 470620 488898
rect 506000 489454 506620 489486
rect 506000 489218 506032 489454
rect 506268 489218 506352 489454
rect 506588 489218 506620 489454
rect 506000 489134 506620 489218
rect 506000 488898 506032 489134
rect 506268 488898 506352 489134
rect 506588 488898 506620 489134
rect 506000 488866 506620 488898
rect 542000 489454 542620 489486
rect 542000 489218 542032 489454
rect 542268 489218 542352 489454
rect 542588 489218 542620 489454
rect 542000 489134 542620 489218
rect 542000 488898 542032 489134
rect 542268 488898 542352 489134
rect 542588 488898 542620 489134
rect 542000 488866 542620 488898
rect 571500 489454 572120 489486
rect 571500 489218 571532 489454
rect 571768 489218 571852 489454
rect 572088 489218 572120 489454
rect 571500 489134 572120 489218
rect 571500 488898 571532 489134
rect 571768 488898 571852 489134
rect 572088 488898 572120 489134
rect 571500 488866 572120 488898
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect 9084 471454 9704 471486
rect 9084 471218 9116 471454
rect 9352 471218 9436 471454
rect 9672 471218 9704 471454
rect 9084 471134 9704 471218
rect 9084 470898 9116 471134
rect 9352 470898 9436 471134
rect 9672 470898 9704 471134
rect 9084 470866 9704 470898
rect 56620 471454 57240 471486
rect 56620 471218 56652 471454
rect 56888 471218 56972 471454
rect 57208 471218 57240 471454
rect 56620 471134 57240 471218
rect 56620 470898 56652 471134
rect 56888 470898 56972 471134
rect 57208 470898 57240 471134
rect 56620 470866 57240 470898
rect 92620 471454 93240 471486
rect 92620 471218 92652 471454
rect 92888 471218 92972 471454
rect 93208 471218 93240 471454
rect 92620 471134 93240 471218
rect 92620 470898 92652 471134
rect 92888 470898 92972 471134
rect 93208 470898 93240 471134
rect 92620 470866 93240 470898
rect 128620 471454 129240 471486
rect 128620 471218 128652 471454
rect 128888 471218 128972 471454
rect 129208 471218 129240 471454
rect 128620 471134 129240 471218
rect 128620 470898 128652 471134
rect 128888 470898 128972 471134
rect 129208 470898 129240 471134
rect 128620 470866 129240 470898
rect 164620 471454 165240 471486
rect 164620 471218 164652 471454
rect 164888 471218 164972 471454
rect 165208 471218 165240 471454
rect 164620 471134 165240 471218
rect 164620 470898 164652 471134
rect 164888 470898 164972 471134
rect 165208 470898 165240 471134
rect 164620 470866 165240 470898
rect 200620 471454 201240 471486
rect 200620 471218 200652 471454
rect 200888 471218 200972 471454
rect 201208 471218 201240 471454
rect 200620 471134 201240 471218
rect 200620 470898 200652 471134
rect 200888 470898 200972 471134
rect 201208 470898 201240 471134
rect 200620 470866 201240 470898
rect 236620 471454 237240 471486
rect 236620 471218 236652 471454
rect 236888 471218 236972 471454
rect 237208 471218 237240 471454
rect 236620 471134 237240 471218
rect 236620 470898 236652 471134
rect 236888 470898 236972 471134
rect 237208 470898 237240 471134
rect 236620 470866 237240 470898
rect 272620 471454 273240 471486
rect 272620 471218 272652 471454
rect 272888 471218 272972 471454
rect 273208 471218 273240 471454
rect 272620 471134 273240 471218
rect 272620 470898 272652 471134
rect 272888 470898 272972 471134
rect 273208 470898 273240 471134
rect 272620 470866 273240 470898
rect 308620 471454 309240 471486
rect 308620 471218 308652 471454
rect 308888 471218 308972 471454
rect 309208 471218 309240 471454
rect 308620 471134 309240 471218
rect 308620 470898 308652 471134
rect 308888 470898 308972 471134
rect 309208 470898 309240 471134
rect 308620 470866 309240 470898
rect 333013 471454 333373 471486
rect 333013 471218 333075 471454
rect 333311 471218 333373 471454
rect 333013 471134 333373 471218
rect 333013 470898 333075 471134
rect 333311 470898 333373 471134
rect 333013 470866 333373 470898
rect 430049 471454 430409 471486
rect 430049 471218 430111 471454
rect 430347 471218 430409 471454
rect 430049 471134 430409 471218
rect 430049 470898 430111 471134
rect 430347 470898 430409 471134
rect 430049 470866 430409 470898
rect 448969 471454 449329 471486
rect 448969 471218 449031 471454
rect 449267 471218 449329 471454
rect 448969 471134 449329 471218
rect 448969 470898 449031 471134
rect 449267 470898 449329 471134
rect 448969 470866 449329 470898
rect 546005 471454 546365 471486
rect 546005 471218 546067 471454
rect 546303 471218 546365 471454
rect 546005 471134 546365 471218
rect 546005 470898 546067 471134
rect 546303 470898 546365 471134
rect 546005 470866 546365 470898
rect 560620 471454 561240 471486
rect 560620 471218 560652 471454
rect 560888 471218 560972 471454
rect 561208 471218 561240 471454
rect 560620 471134 561240 471218
rect 560620 470898 560652 471134
rect 560888 470898 560972 471134
rect 561208 470898 561240 471134
rect 560620 470866 561240 470898
rect 570260 471454 570880 471486
rect 570260 471218 570292 471454
rect 570528 471218 570612 471454
rect 570848 471218 570880 471454
rect 570260 471134 570880 471218
rect 570260 470898 570292 471134
rect 570528 470898 570612 471134
rect 570848 470898 570880 471134
rect 570260 470866 570880 470898
rect 7844 453454 8464 453486
rect 7844 453218 7876 453454
rect 8112 453218 8196 453454
rect 8432 453218 8464 453454
rect 7844 453134 8464 453218
rect 7844 452898 7876 453134
rect 8112 452898 8196 453134
rect 8432 452898 8464 453134
rect 7844 452866 8464 452898
rect 38000 453454 38620 453486
rect 38000 453218 38032 453454
rect 38268 453218 38352 453454
rect 38588 453218 38620 453454
rect 38000 453134 38620 453218
rect 38000 452898 38032 453134
rect 38268 452898 38352 453134
rect 38588 452898 38620 453134
rect 38000 452866 38620 452898
rect 74000 453454 74620 453486
rect 74000 453218 74032 453454
rect 74268 453218 74352 453454
rect 74588 453218 74620 453454
rect 74000 453134 74620 453218
rect 74000 452898 74032 453134
rect 74268 452898 74352 453134
rect 74588 452898 74620 453134
rect 74000 452866 74620 452898
rect 110000 453454 110620 453486
rect 110000 453218 110032 453454
rect 110268 453218 110352 453454
rect 110588 453218 110620 453454
rect 110000 453134 110620 453218
rect 110000 452898 110032 453134
rect 110268 452898 110352 453134
rect 110588 452898 110620 453134
rect 110000 452866 110620 452898
rect 146000 453454 146620 453486
rect 146000 453218 146032 453454
rect 146268 453218 146352 453454
rect 146588 453218 146620 453454
rect 146000 453134 146620 453218
rect 146000 452898 146032 453134
rect 146268 452898 146352 453134
rect 146588 452898 146620 453134
rect 146000 452866 146620 452898
rect 182000 453454 182620 453486
rect 182000 453218 182032 453454
rect 182268 453218 182352 453454
rect 182588 453218 182620 453454
rect 182000 453134 182620 453218
rect 182000 452898 182032 453134
rect 182268 452898 182352 453134
rect 182588 452898 182620 453134
rect 182000 452866 182620 452898
rect 218000 453454 218620 453486
rect 218000 453218 218032 453454
rect 218268 453218 218352 453454
rect 218588 453218 218620 453454
rect 218000 453134 218620 453218
rect 218000 452898 218032 453134
rect 218268 452898 218352 453134
rect 218588 452898 218620 453134
rect 218000 452866 218620 452898
rect 254000 453454 254620 453486
rect 254000 453218 254032 453454
rect 254268 453218 254352 453454
rect 254588 453218 254620 453454
rect 254000 453134 254620 453218
rect 254000 452898 254032 453134
rect 254268 452898 254352 453134
rect 254588 452898 254620 453134
rect 254000 452866 254620 452898
rect 290000 453454 290620 453486
rect 290000 453218 290032 453454
rect 290268 453218 290352 453454
rect 290588 453218 290620 453454
rect 290000 453134 290620 453218
rect 290000 452898 290032 453134
rect 290268 452898 290352 453134
rect 290588 452898 290620 453134
rect 290000 452866 290620 452898
rect 326000 453454 326620 453486
rect 326000 453218 326032 453454
rect 326268 453218 326352 453454
rect 326588 453218 326620 453454
rect 326000 453134 326620 453218
rect 326000 452898 326032 453134
rect 326268 452898 326352 453134
rect 326588 452898 326620 453134
rect 326000 452866 326620 452898
rect 332293 453454 332653 453486
rect 332293 453218 332355 453454
rect 332591 453218 332653 453454
rect 332293 453134 332653 453218
rect 332293 452898 332355 453134
rect 332591 452898 332653 453134
rect 332293 452866 332653 452898
rect 430769 453454 431129 453486
rect 430769 453218 430831 453454
rect 431067 453218 431129 453454
rect 430769 453134 431129 453218
rect 430769 452898 430831 453134
rect 431067 452898 431129 453134
rect 430769 452866 431129 452898
rect 434000 453454 434620 453486
rect 434000 453218 434032 453454
rect 434268 453218 434352 453454
rect 434588 453218 434620 453454
rect 434000 453134 434620 453218
rect 434000 452898 434032 453134
rect 434268 452898 434352 453134
rect 434588 452898 434620 453134
rect 434000 452866 434620 452898
rect 448249 453454 448609 453486
rect 448249 453218 448311 453454
rect 448547 453218 448609 453454
rect 448249 453134 448609 453218
rect 448249 452898 448311 453134
rect 448547 452898 448609 453134
rect 448249 452866 448609 452898
rect 546725 453454 547085 453486
rect 546725 453218 546787 453454
rect 547023 453218 547085 453454
rect 546725 453134 547085 453218
rect 546725 452898 546787 453134
rect 547023 452898 547085 453134
rect 546725 452866 547085 452898
rect 571500 453454 572120 453486
rect 571500 453218 571532 453454
rect 571768 453218 571852 453454
rect 572088 453218 572120 453454
rect 571500 453134 572120 453218
rect 571500 452898 571532 453134
rect 571768 452898 571852 453134
rect 572088 452898 572120 453134
rect 571500 452866 572120 452898
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect 9084 435454 9704 435486
rect 9084 435218 9116 435454
rect 9352 435218 9436 435454
rect 9672 435218 9704 435454
rect 9084 435134 9704 435218
rect 9084 434898 9116 435134
rect 9352 434898 9436 435134
rect 9672 434898 9704 435134
rect 9084 434866 9704 434898
rect 56620 435454 57240 435486
rect 56620 435218 56652 435454
rect 56888 435218 56972 435454
rect 57208 435218 57240 435454
rect 56620 435134 57240 435218
rect 56620 434898 56652 435134
rect 56888 434898 56972 435134
rect 57208 434898 57240 435134
rect 56620 434866 57240 434898
rect 92620 435454 93240 435486
rect 92620 435218 92652 435454
rect 92888 435218 92972 435454
rect 93208 435218 93240 435454
rect 92620 435134 93240 435218
rect 92620 434898 92652 435134
rect 92888 434898 92972 435134
rect 93208 434898 93240 435134
rect 92620 434866 93240 434898
rect 128620 435454 129240 435486
rect 128620 435218 128652 435454
rect 128888 435218 128972 435454
rect 129208 435218 129240 435454
rect 128620 435134 129240 435218
rect 128620 434898 128652 435134
rect 128888 434898 128972 435134
rect 129208 434898 129240 435134
rect 128620 434866 129240 434898
rect 164620 435454 165240 435486
rect 164620 435218 164652 435454
rect 164888 435218 164972 435454
rect 165208 435218 165240 435454
rect 164620 435134 165240 435218
rect 164620 434898 164652 435134
rect 164888 434898 164972 435134
rect 165208 434898 165240 435134
rect 164620 434866 165240 434898
rect 200620 435454 201240 435486
rect 200620 435218 200652 435454
rect 200888 435218 200972 435454
rect 201208 435218 201240 435454
rect 200620 435134 201240 435218
rect 200620 434898 200652 435134
rect 200888 434898 200972 435134
rect 201208 434898 201240 435134
rect 200620 434866 201240 434898
rect 236620 435454 237240 435486
rect 236620 435218 236652 435454
rect 236888 435218 236972 435454
rect 237208 435218 237240 435454
rect 236620 435134 237240 435218
rect 236620 434898 236652 435134
rect 236888 434898 236972 435134
rect 237208 434898 237240 435134
rect 236620 434866 237240 434898
rect 272620 435454 273240 435486
rect 272620 435218 272652 435454
rect 272888 435218 272972 435454
rect 273208 435218 273240 435454
rect 272620 435134 273240 435218
rect 272620 434898 272652 435134
rect 272888 434898 272972 435134
rect 273208 434898 273240 435134
rect 272620 434866 273240 434898
rect 308620 435454 309240 435486
rect 308620 435218 308652 435454
rect 308888 435218 308972 435454
rect 309208 435218 309240 435454
rect 308620 435134 309240 435218
rect 308620 434898 308652 435134
rect 308888 434898 308972 435134
rect 309208 434898 309240 435134
rect 308620 434866 309240 434898
rect 333013 435454 333373 435486
rect 333013 435218 333075 435454
rect 333311 435218 333373 435454
rect 333013 435134 333373 435218
rect 333013 434898 333075 435134
rect 333311 434898 333373 435134
rect 333013 434866 333373 434898
rect 430049 435454 430409 435486
rect 430049 435218 430111 435454
rect 430347 435218 430409 435454
rect 430049 435134 430409 435218
rect 430049 434898 430111 435134
rect 430347 434898 430409 435134
rect 430049 434866 430409 434898
rect 448969 435454 449329 435486
rect 448969 435218 449031 435454
rect 449267 435218 449329 435454
rect 448969 435134 449329 435218
rect 448969 434898 449031 435134
rect 449267 434898 449329 435134
rect 448969 434866 449329 434898
rect 546005 435454 546365 435486
rect 546005 435218 546067 435454
rect 546303 435218 546365 435454
rect 546005 435134 546365 435218
rect 546005 434898 546067 435134
rect 546303 434898 546365 435134
rect 546005 434866 546365 434898
rect 560620 435454 561240 435486
rect 560620 435218 560652 435454
rect 560888 435218 560972 435454
rect 561208 435218 561240 435454
rect 560620 435134 561240 435218
rect 560620 434898 560652 435134
rect 560888 434898 560972 435134
rect 561208 434898 561240 435134
rect 560620 434866 561240 434898
rect 570260 435454 570880 435486
rect 570260 435218 570292 435454
rect 570528 435218 570612 435454
rect 570848 435218 570880 435454
rect 570260 435134 570880 435218
rect 570260 434898 570292 435134
rect 570528 434898 570612 435134
rect 570848 434898 570880 435134
rect 570260 434866 570880 434898
rect 7844 417454 8464 417486
rect 7844 417218 7876 417454
rect 8112 417218 8196 417454
rect 8432 417218 8464 417454
rect 7844 417134 8464 417218
rect 7844 416898 7876 417134
rect 8112 416898 8196 417134
rect 8432 416898 8464 417134
rect 7844 416866 8464 416898
rect 38000 417454 38620 417486
rect 38000 417218 38032 417454
rect 38268 417218 38352 417454
rect 38588 417218 38620 417454
rect 38000 417134 38620 417218
rect 38000 416898 38032 417134
rect 38268 416898 38352 417134
rect 38588 416898 38620 417134
rect 38000 416866 38620 416898
rect 74000 417454 74620 417486
rect 74000 417218 74032 417454
rect 74268 417218 74352 417454
rect 74588 417218 74620 417454
rect 74000 417134 74620 417218
rect 74000 416898 74032 417134
rect 74268 416898 74352 417134
rect 74588 416898 74620 417134
rect 74000 416866 74620 416898
rect 110000 417454 110620 417486
rect 110000 417218 110032 417454
rect 110268 417218 110352 417454
rect 110588 417218 110620 417454
rect 110000 417134 110620 417218
rect 110000 416898 110032 417134
rect 110268 416898 110352 417134
rect 110588 416898 110620 417134
rect 110000 416866 110620 416898
rect 146000 417454 146620 417486
rect 146000 417218 146032 417454
rect 146268 417218 146352 417454
rect 146588 417218 146620 417454
rect 146000 417134 146620 417218
rect 146000 416898 146032 417134
rect 146268 416898 146352 417134
rect 146588 416898 146620 417134
rect 146000 416866 146620 416898
rect 182000 417454 182620 417486
rect 182000 417218 182032 417454
rect 182268 417218 182352 417454
rect 182588 417218 182620 417454
rect 182000 417134 182620 417218
rect 182000 416898 182032 417134
rect 182268 416898 182352 417134
rect 182588 416898 182620 417134
rect 182000 416866 182620 416898
rect 218000 417454 218620 417486
rect 218000 417218 218032 417454
rect 218268 417218 218352 417454
rect 218588 417218 218620 417454
rect 218000 417134 218620 417218
rect 218000 416898 218032 417134
rect 218268 416898 218352 417134
rect 218588 416898 218620 417134
rect 218000 416866 218620 416898
rect 254000 417454 254620 417486
rect 254000 417218 254032 417454
rect 254268 417218 254352 417454
rect 254588 417218 254620 417454
rect 254000 417134 254620 417218
rect 254000 416898 254032 417134
rect 254268 416898 254352 417134
rect 254588 416898 254620 417134
rect 254000 416866 254620 416898
rect 290000 417454 290620 417486
rect 290000 417218 290032 417454
rect 290268 417218 290352 417454
rect 290588 417218 290620 417454
rect 290000 417134 290620 417218
rect 290000 416898 290032 417134
rect 290268 416898 290352 417134
rect 290588 416898 290620 417134
rect 290000 416866 290620 416898
rect 326000 417454 326620 417486
rect 326000 417218 326032 417454
rect 326268 417218 326352 417454
rect 326588 417218 326620 417454
rect 326000 417134 326620 417218
rect 326000 416898 326032 417134
rect 326268 416898 326352 417134
rect 326588 416898 326620 417134
rect 326000 416866 326620 416898
rect 332293 417454 332653 417486
rect 332293 417218 332355 417454
rect 332591 417218 332653 417454
rect 332293 417134 332653 417218
rect 332293 416898 332355 417134
rect 332591 416898 332653 417134
rect 332293 416866 332653 416898
rect 430769 417454 431129 417486
rect 430769 417218 430831 417454
rect 431067 417218 431129 417454
rect 430769 417134 431129 417218
rect 430769 416898 430831 417134
rect 431067 416898 431129 417134
rect 430769 416866 431129 416898
rect 434000 417454 434620 417486
rect 434000 417218 434032 417454
rect 434268 417218 434352 417454
rect 434588 417218 434620 417454
rect 434000 417134 434620 417218
rect 434000 416898 434032 417134
rect 434268 416898 434352 417134
rect 434588 416898 434620 417134
rect 434000 416866 434620 416898
rect 448249 417454 448609 417486
rect 448249 417218 448311 417454
rect 448547 417218 448609 417454
rect 448249 417134 448609 417218
rect 448249 416898 448311 417134
rect 448547 416898 448609 417134
rect 448249 416866 448609 416898
rect 546725 417454 547085 417486
rect 546725 417218 546787 417454
rect 547023 417218 547085 417454
rect 546725 417134 547085 417218
rect 546725 416898 546787 417134
rect 547023 416898 547085 417134
rect 546725 416866 547085 416898
rect 571500 417454 572120 417486
rect 571500 417218 571532 417454
rect 571768 417218 571852 417454
rect 572088 417218 572120 417454
rect 571500 417134 572120 417218
rect 571500 416898 571532 417134
rect 571768 416898 571852 417134
rect 572088 416898 572120 417134
rect 571500 416866 572120 416898
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect 9084 399454 9704 399486
rect 9084 399218 9116 399454
rect 9352 399218 9436 399454
rect 9672 399218 9704 399454
rect 9084 399134 9704 399218
rect 9084 398898 9116 399134
rect 9352 398898 9436 399134
rect 9672 398898 9704 399134
rect 9084 398866 9704 398898
rect 56620 399454 57240 399486
rect 56620 399218 56652 399454
rect 56888 399218 56972 399454
rect 57208 399218 57240 399454
rect 56620 399134 57240 399218
rect 56620 398898 56652 399134
rect 56888 398898 56972 399134
rect 57208 398898 57240 399134
rect 56620 398866 57240 398898
rect 92620 399454 93240 399486
rect 92620 399218 92652 399454
rect 92888 399218 92972 399454
rect 93208 399218 93240 399454
rect 92620 399134 93240 399218
rect 92620 398898 92652 399134
rect 92888 398898 92972 399134
rect 93208 398898 93240 399134
rect 92620 398866 93240 398898
rect 128620 399454 129240 399486
rect 128620 399218 128652 399454
rect 128888 399218 128972 399454
rect 129208 399218 129240 399454
rect 128620 399134 129240 399218
rect 128620 398898 128652 399134
rect 128888 398898 128972 399134
rect 129208 398898 129240 399134
rect 128620 398866 129240 398898
rect 164620 399454 165240 399486
rect 164620 399218 164652 399454
rect 164888 399218 164972 399454
rect 165208 399218 165240 399454
rect 164620 399134 165240 399218
rect 164620 398898 164652 399134
rect 164888 398898 164972 399134
rect 165208 398898 165240 399134
rect 164620 398866 165240 398898
rect 200620 399454 201240 399486
rect 200620 399218 200652 399454
rect 200888 399218 200972 399454
rect 201208 399218 201240 399454
rect 200620 399134 201240 399218
rect 200620 398898 200652 399134
rect 200888 398898 200972 399134
rect 201208 398898 201240 399134
rect 200620 398866 201240 398898
rect 236620 399454 237240 399486
rect 236620 399218 236652 399454
rect 236888 399218 236972 399454
rect 237208 399218 237240 399454
rect 236620 399134 237240 399218
rect 236620 398898 236652 399134
rect 236888 398898 236972 399134
rect 237208 398898 237240 399134
rect 236620 398866 237240 398898
rect 272620 399454 273240 399486
rect 272620 399218 272652 399454
rect 272888 399218 272972 399454
rect 273208 399218 273240 399454
rect 272620 399134 273240 399218
rect 272620 398898 272652 399134
rect 272888 398898 272972 399134
rect 273208 398898 273240 399134
rect 272620 398866 273240 398898
rect 308620 399454 309240 399486
rect 308620 399218 308652 399454
rect 308888 399218 308972 399454
rect 309208 399218 309240 399454
rect 308620 399134 309240 399218
rect 308620 398898 308652 399134
rect 308888 398898 308972 399134
rect 309208 398898 309240 399134
rect 308620 398866 309240 398898
rect 333013 399454 333373 399486
rect 333013 399218 333075 399454
rect 333311 399218 333373 399454
rect 333013 399134 333373 399218
rect 333013 398898 333075 399134
rect 333311 398898 333373 399134
rect 333013 398866 333373 398898
rect 430049 399454 430409 399486
rect 430049 399218 430111 399454
rect 430347 399218 430409 399454
rect 430049 399134 430409 399218
rect 430049 398898 430111 399134
rect 430347 398898 430409 399134
rect 430049 398866 430409 398898
rect 448969 399454 449329 399486
rect 448969 399218 449031 399454
rect 449267 399218 449329 399454
rect 448969 399134 449329 399218
rect 448969 398898 449031 399134
rect 449267 398898 449329 399134
rect 448969 398866 449329 398898
rect 546005 399454 546365 399486
rect 546005 399218 546067 399454
rect 546303 399218 546365 399454
rect 546005 399134 546365 399218
rect 546005 398898 546067 399134
rect 546303 398898 546365 399134
rect 546005 398866 546365 398898
rect 560620 399454 561240 399486
rect 560620 399218 560652 399454
rect 560888 399218 560972 399454
rect 561208 399218 561240 399454
rect 560620 399134 561240 399218
rect 560620 398898 560652 399134
rect 560888 398898 560972 399134
rect 561208 398898 561240 399134
rect 560620 398866 561240 398898
rect 570260 399454 570880 399486
rect 570260 399218 570292 399454
rect 570528 399218 570612 399454
rect 570848 399218 570880 399454
rect 570260 399134 570880 399218
rect 570260 398898 570292 399134
rect 570528 398898 570612 399134
rect 570848 398898 570880 399134
rect 570260 398866 570880 398898
rect 7844 381454 8464 381486
rect 7844 381218 7876 381454
rect 8112 381218 8196 381454
rect 8432 381218 8464 381454
rect 7844 381134 8464 381218
rect 7844 380898 7876 381134
rect 8112 380898 8196 381134
rect 8432 380898 8464 381134
rect 7844 380866 8464 380898
rect 38000 381454 38620 381486
rect 38000 381218 38032 381454
rect 38268 381218 38352 381454
rect 38588 381218 38620 381454
rect 38000 381134 38620 381218
rect 38000 380898 38032 381134
rect 38268 380898 38352 381134
rect 38588 380898 38620 381134
rect 38000 380866 38620 380898
rect 74000 381454 74620 381486
rect 74000 381218 74032 381454
rect 74268 381218 74352 381454
rect 74588 381218 74620 381454
rect 74000 381134 74620 381218
rect 74000 380898 74032 381134
rect 74268 380898 74352 381134
rect 74588 380898 74620 381134
rect 74000 380866 74620 380898
rect 110000 381454 110620 381486
rect 110000 381218 110032 381454
rect 110268 381218 110352 381454
rect 110588 381218 110620 381454
rect 110000 381134 110620 381218
rect 110000 380898 110032 381134
rect 110268 380898 110352 381134
rect 110588 380898 110620 381134
rect 110000 380866 110620 380898
rect 146000 381454 146620 381486
rect 146000 381218 146032 381454
rect 146268 381218 146352 381454
rect 146588 381218 146620 381454
rect 146000 381134 146620 381218
rect 146000 380898 146032 381134
rect 146268 380898 146352 381134
rect 146588 380898 146620 381134
rect 146000 380866 146620 380898
rect 182000 381454 182620 381486
rect 182000 381218 182032 381454
rect 182268 381218 182352 381454
rect 182588 381218 182620 381454
rect 182000 381134 182620 381218
rect 182000 380898 182032 381134
rect 182268 380898 182352 381134
rect 182588 380898 182620 381134
rect 182000 380866 182620 380898
rect 218000 381454 218620 381486
rect 218000 381218 218032 381454
rect 218268 381218 218352 381454
rect 218588 381218 218620 381454
rect 218000 381134 218620 381218
rect 218000 380898 218032 381134
rect 218268 380898 218352 381134
rect 218588 380898 218620 381134
rect 218000 380866 218620 380898
rect 254000 381454 254620 381486
rect 254000 381218 254032 381454
rect 254268 381218 254352 381454
rect 254588 381218 254620 381454
rect 254000 381134 254620 381218
rect 254000 380898 254032 381134
rect 254268 380898 254352 381134
rect 254588 380898 254620 381134
rect 254000 380866 254620 380898
rect 290000 381454 290620 381486
rect 290000 381218 290032 381454
rect 290268 381218 290352 381454
rect 290588 381218 290620 381454
rect 290000 381134 290620 381218
rect 290000 380898 290032 381134
rect 290268 380898 290352 381134
rect 290588 380898 290620 381134
rect 290000 380866 290620 380898
rect 326000 381454 326620 381486
rect 326000 381218 326032 381454
rect 326268 381218 326352 381454
rect 326588 381218 326620 381454
rect 326000 381134 326620 381218
rect 326000 380898 326032 381134
rect 326268 380898 326352 381134
rect 326588 380898 326620 381134
rect 326000 380866 326620 380898
rect 362000 381454 362620 381486
rect 362000 381218 362032 381454
rect 362268 381218 362352 381454
rect 362588 381218 362620 381454
rect 362000 381134 362620 381218
rect 362000 380898 362032 381134
rect 362268 380898 362352 381134
rect 362588 380898 362620 381134
rect 362000 380866 362620 380898
rect 398000 381454 398620 381486
rect 398000 381218 398032 381454
rect 398268 381218 398352 381454
rect 398588 381218 398620 381454
rect 398000 381134 398620 381218
rect 398000 380898 398032 381134
rect 398268 380898 398352 381134
rect 398588 380898 398620 381134
rect 398000 380866 398620 380898
rect 434000 381454 434620 381486
rect 434000 381218 434032 381454
rect 434268 381218 434352 381454
rect 434588 381218 434620 381454
rect 434000 381134 434620 381218
rect 434000 380898 434032 381134
rect 434268 380898 434352 381134
rect 434588 380898 434620 381134
rect 434000 380866 434620 380898
rect 470000 381454 470620 381486
rect 470000 381218 470032 381454
rect 470268 381218 470352 381454
rect 470588 381218 470620 381454
rect 470000 381134 470620 381218
rect 470000 380898 470032 381134
rect 470268 380898 470352 381134
rect 470588 380898 470620 381134
rect 470000 380866 470620 380898
rect 506000 381454 506620 381486
rect 506000 381218 506032 381454
rect 506268 381218 506352 381454
rect 506588 381218 506620 381454
rect 506000 381134 506620 381218
rect 506000 380898 506032 381134
rect 506268 380898 506352 381134
rect 506588 380898 506620 381134
rect 506000 380866 506620 380898
rect 542000 381454 542620 381486
rect 542000 381218 542032 381454
rect 542268 381218 542352 381454
rect 542588 381218 542620 381454
rect 542000 381134 542620 381218
rect 542000 380898 542032 381134
rect 542268 380898 542352 381134
rect 542588 380898 542620 381134
rect 542000 380866 542620 380898
rect 571500 381454 572120 381486
rect 571500 381218 571532 381454
rect 571768 381218 571852 381454
rect 572088 381218 572120 381454
rect 571500 381134 572120 381218
rect 571500 380898 571532 381134
rect 571768 380898 571852 381134
rect 572088 380898 572120 381134
rect 571500 380866 572120 380898
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect 9084 363454 9704 363486
rect 9084 363218 9116 363454
rect 9352 363218 9436 363454
rect 9672 363218 9704 363454
rect 9084 363134 9704 363218
rect 9084 362898 9116 363134
rect 9352 362898 9436 363134
rect 9672 362898 9704 363134
rect 9084 362866 9704 362898
rect 56620 363454 57240 363486
rect 56620 363218 56652 363454
rect 56888 363218 56972 363454
rect 57208 363218 57240 363454
rect 56620 363134 57240 363218
rect 56620 362898 56652 363134
rect 56888 362898 56972 363134
rect 57208 362898 57240 363134
rect 56620 362866 57240 362898
rect 92620 363454 93240 363486
rect 92620 363218 92652 363454
rect 92888 363218 92972 363454
rect 93208 363218 93240 363454
rect 92620 363134 93240 363218
rect 92620 362898 92652 363134
rect 92888 362898 92972 363134
rect 93208 362898 93240 363134
rect 92620 362866 93240 362898
rect 128620 363454 129240 363486
rect 128620 363218 128652 363454
rect 128888 363218 128972 363454
rect 129208 363218 129240 363454
rect 128620 363134 129240 363218
rect 128620 362898 128652 363134
rect 128888 362898 128972 363134
rect 129208 362898 129240 363134
rect 128620 362866 129240 362898
rect 164620 363454 165240 363486
rect 164620 363218 164652 363454
rect 164888 363218 164972 363454
rect 165208 363218 165240 363454
rect 164620 363134 165240 363218
rect 164620 362898 164652 363134
rect 164888 362898 164972 363134
rect 165208 362898 165240 363134
rect 164620 362866 165240 362898
rect 200620 363454 201240 363486
rect 200620 363218 200652 363454
rect 200888 363218 200972 363454
rect 201208 363218 201240 363454
rect 200620 363134 201240 363218
rect 200620 362898 200652 363134
rect 200888 362898 200972 363134
rect 201208 362898 201240 363134
rect 200620 362866 201240 362898
rect 236620 363454 237240 363486
rect 236620 363218 236652 363454
rect 236888 363218 236972 363454
rect 237208 363218 237240 363454
rect 236620 363134 237240 363218
rect 236620 362898 236652 363134
rect 236888 362898 236972 363134
rect 237208 362898 237240 363134
rect 236620 362866 237240 362898
rect 272620 363454 273240 363486
rect 272620 363218 272652 363454
rect 272888 363218 272972 363454
rect 273208 363218 273240 363454
rect 272620 363134 273240 363218
rect 272620 362898 272652 363134
rect 272888 362898 272972 363134
rect 273208 362898 273240 363134
rect 272620 362866 273240 362898
rect 308620 363454 309240 363486
rect 308620 363218 308652 363454
rect 308888 363218 308972 363454
rect 309208 363218 309240 363454
rect 308620 363134 309240 363218
rect 308620 362898 308652 363134
rect 308888 362898 308972 363134
rect 309208 362898 309240 363134
rect 308620 362866 309240 362898
rect 333013 363454 333373 363486
rect 333013 363218 333075 363454
rect 333311 363218 333373 363454
rect 333013 363134 333373 363218
rect 333013 362898 333075 363134
rect 333311 362898 333373 363134
rect 333013 362866 333373 362898
rect 430049 363454 430409 363486
rect 430049 363218 430111 363454
rect 430347 363218 430409 363454
rect 430049 363134 430409 363218
rect 430049 362898 430111 363134
rect 430347 362898 430409 363134
rect 430049 362866 430409 362898
rect 448969 363454 449329 363486
rect 448969 363218 449031 363454
rect 449267 363218 449329 363454
rect 448969 363134 449329 363218
rect 448969 362898 449031 363134
rect 449267 362898 449329 363134
rect 448969 362866 449329 362898
rect 546005 363454 546365 363486
rect 546005 363218 546067 363454
rect 546303 363218 546365 363454
rect 546005 363134 546365 363218
rect 546005 362898 546067 363134
rect 546303 362898 546365 363134
rect 546005 362866 546365 362898
rect 560620 363454 561240 363486
rect 560620 363218 560652 363454
rect 560888 363218 560972 363454
rect 561208 363218 561240 363454
rect 560620 363134 561240 363218
rect 560620 362898 560652 363134
rect 560888 362898 560972 363134
rect 561208 362898 561240 363134
rect 560620 362866 561240 362898
rect 570260 363454 570880 363486
rect 570260 363218 570292 363454
rect 570528 363218 570612 363454
rect 570848 363218 570880 363454
rect 570260 363134 570880 363218
rect 570260 362898 570292 363134
rect 570528 362898 570612 363134
rect 570848 362898 570880 363134
rect 570260 362866 570880 362898
rect 7844 345454 8464 345486
rect 7844 345218 7876 345454
rect 8112 345218 8196 345454
rect 8432 345218 8464 345454
rect 7844 345134 8464 345218
rect 7844 344898 7876 345134
rect 8112 344898 8196 345134
rect 8432 344898 8464 345134
rect 7844 344866 8464 344898
rect 38000 345454 38620 345486
rect 38000 345218 38032 345454
rect 38268 345218 38352 345454
rect 38588 345218 38620 345454
rect 38000 345134 38620 345218
rect 38000 344898 38032 345134
rect 38268 344898 38352 345134
rect 38588 344898 38620 345134
rect 38000 344866 38620 344898
rect 74000 345454 74620 345486
rect 74000 345218 74032 345454
rect 74268 345218 74352 345454
rect 74588 345218 74620 345454
rect 74000 345134 74620 345218
rect 74000 344898 74032 345134
rect 74268 344898 74352 345134
rect 74588 344898 74620 345134
rect 74000 344866 74620 344898
rect 110000 345454 110620 345486
rect 110000 345218 110032 345454
rect 110268 345218 110352 345454
rect 110588 345218 110620 345454
rect 110000 345134 110620 345218
rect 110000 344898 110032 345134
rect 110268 344898 110352 345134
rect 110588 344898 110620 345134
rect 110000 344866 110620 344898
rect 146000 345454 146620 345486
rect 146000 345218 146032 345454
rect 146268 345218 146352 345454
rect 146588 345218 146620 345454
rect 146000 345134 146620 345218
rect 146000 344898 146032 345134
rect 146268 344898 146352 345134
rect 146588 344898 146620 345134
rect 146000 344866 146620 344898
rect 182000 345454 182620 345486
rect 182000 345218 182032 345454
rect 182268 345218 182352 345454
rect 182588 345218 182620 345454
rect 182000 345134 182620 345218
rect 182000 344898 182032 345134
rect 182268 344898 182352 345134
rect 182588 344898 182620 345134
rect 182000 344866 182620 344898
rect 218000 345454 218620 345486
rect 218000 345218 218032 345454
rect 218268 345218 218352 345454
rect 218588 345218 218620 345454
rect 218000 345134 218620 345218
rect 218000 344898 218032 345134
rect 218268 344898 218352 345134
rect 218588 344898 218620 345134
rect 218000 344866 218620 344898
rect 254000 345454 254620 345486
rect 254000 345218 254032 345454
rect 254268 345218 254352 345454
rect 254588 345218 254620 345454
rect 254000 345134 254620 345218
rect 254000 344898 254032 345134
rect 254268 344898 254352 345134
rect 254588 344898 254620 345134
rect 254000 344866 254620 344898
rect 290000 345454 290620 345486
rect 290000 345218 290032 345454
rect 290268 345218 290352 345454
rect 290588 345218 290620 345454
rect 290000 345134 290620 345218
rect 290000 344898 290032 345134
rect 290268 344898 290352 345134
rect 290588 344898 290620 345134
rect 290000 344866 290620 344898
rect 326000 345454 326620 345486
rect 326000 345218 326032 345454
rect 326268 345218 326352 345454
rect 326588 345218 326620 345454
rect 326000 345134 326620 345218
rect 326000 344898 326032 345134
rect 326268 344898 326352 345134
rect 326588 344898 326620 345134
rect 326000 344866 326620 344898
rect 332293 345454 332653 345486
rect 332293 345218 332355 345454
rect 332591 345218 332653 345454
rect 332293 345134 332653 345218
rect 332293 344898 332355 345134
rect 332591 344898 332653 345134
rect 332293 344866 332653 344898
rect 430769 345454 431129 345486
rect 430769 345218 430831 345454
rect 431067 345218 431129 345454
rect 430769 345134 431129 345218
rect 430769 344898 430831 345134
rect 431067 344898 431129 345134
rect 430769 344866 431129 344898
rect 434000 345454 434620 345486
rect 434000 345218 434032 345454
rect 434268 345218 434352 345454
rect 434588 345218 434620 345454
rect 434000 345134 434620 345218
rect 434000 344898 434032 345134
rect 434268 344898 434352 345134
rect 434588 344898 434620 345134
rect 434000 344866 434620 344898
rect 448249 345454 448609 345486
rect 448249 345218 448311 345454
rect 448547 345218 448609 345454
rect 448249 345134 448609 345218
rect 448249 344898 448311 345134
rect 448547 344898 448609 345134
rect 448249 344866 448609 344898
rect 546725 345454 547085 345486
rect 546725 345218 546787 345454
rect 547023 345218 547085 345454
rect 546725 345134 547085 345218
rect 546725 344898 546787 345134
rect 547023 344898 547085 345134
rect 546725 344866 547085 344898
rect 571500 345454 572120 345486
rect 571500 345218 571532 345454
rect 571768 345218 571852 345454
rect 572088 345218 572120 345454
rect 571500 345134 572120 345218
rect 571500 344898 571532 345134
rect 571768 344898 571852 345134
rect 572088 344898 572120 345134
rect 571500 344866 572120 344898
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect 9084 327454 9704 327486
rect 9084 327218 9116 327454
rect 9352 327218 9436 327454
rect 9672 327218 9704 327454
rect 9084 327134 9704 327218
rect 9084 326898 9116 327134
rect 9352 326898 9436 327134
rect 9672 326898 9704 327134
rect 9084 326866 9704 326898
rect 56620 327454 57240 327486
rect 56620 327218 56652 327454
rect 56888 327218 56972 327454
rect 57208 327218 57240 327454
rect 56620 327134 57240 327218
rect 56620 326898 56652 327134
rect 56888 326898 56972 327134
rect 57208 326898 57240 327134
rect 56620 326866 57240 326898
rect 92620 327454 93240 327486
rect 92620 327218 92652 327454
rect 92888 327218 92972 327454
rect 93208 327218 93240 327454
rect 92620 327134 93240 327218
rect 92620 326898 92652 327134
rect 92888 326898 92972 327134
rect 93208 326898 93240 327134
rect 92620 326866 93240 326898
rect 128620 327454 129240 327486
rect 128620 327218 128652 327454
rect 128888 327218 128972 327454
rect 129208 327218 129240 327454
rect 128620 327134 129240 327218
rect 128620 326898 128652 327134
rect 128888 326898 128972 327134
rect 129208 326898 129240 327134
rect 128620 326866 129240 326898
rect 164620 327454 165240 327486
rect 164620 327218 164652 327454
rect 164888 327218 164972 327454
rect 165208 327218 165240 327454
rect 164620 327134 165240 327218
rect 164620 326898 164652 327134
rect 164888 326898 164972 327134
rect 165208 326898 165240 327134
rect 164620 326866 165240 326898
rect 200620 327454 201240 327486
rect 200620 327218 200652 327454
rect 200888 327218 200972 327454
rect 201208 327218 201240 327454
rect 200620 327134 201240 327218
rect 200620 326898 200652 327134
rect 200888 326898 200972 327134
rect 201208 326898 201240 327134
rect 200620 326866 201240 326898
rect 236620 327454 237240 327486
rect 236620 327218 236652 327454
rect 236888 327218 236972 327454
rect 237208 327218 237240 327454
rect 236620 327134 237240 327218
rect 236620 326898 236652 327134
rect 236888 326898 236972 327134
rect 237208 326898 237240 327134
rect 236620 326866 237240 326898
rect 272620 327454 273240 327486
rect 272620 327218 272652 327454
rect 272888 327218 272972 327454
rect 273208 327218 273240 327454
rect 272620 327134 273240 327218
rect 272620 326898 272652 327134
rect 272888 326898 272972 327134
rect 273208 326898 273240 327134
rect 272620 326866 273240 326898
rect 308620 327454 309240 327486
rect 308620 327218 308652 327454
rect 308888 327218 308972 327454
rect 309208 327218 309240 327454
rect 308620 327134 309240 327218
rect 308620 326898 308652 327134
rect 308888 326898 308972 327134
rect 309208 326898 309240 327134
rect 308620 326866 309240 326898
rect 333013 327454 333373 327486
rect 333013 327218 333075 327454
rect 333311 327218 333373 327454
rect 333013 327134 333373 327218
rect 333013 326898 333075 327134
rect 333311 326898 333373 327134
rect 333013 326866 333373 326898
rect 430049 327454 430409 327486
rect 430049 327218 430111 327454
rect 430347 327218 430409 327454
rect 430049 327134 430409 327218
rect 430049 326898 430111 327134
rect 430347 326898 430409 327134
rect 430049 326866 430409 326898
rect 448969 327454 449329 327486
rect 448969 327218 449031 327454
rect 449267 327218 449329 327454
rect 448969 327134 449329 327218
rect 448969 326898 449031 327134
rect 449267 326898 449329 327134
rect 448969 326866 449329 326898
rect 546005 327454 546365 327486
rect 546005 327218 546067 327454
rect 546303 327218 546365 327454
rect 546005 327134 546365 327218
rect 546005 326898 546067 327134
rect 546303 326898 546365 327134
rect 546005 326866 546365 326898
rect 560620 327454 561240 327486
rect 560620 327218 560652 327454
rect 560888 327218 560972 327454
rect 561208 327218 561240 327454
rect 560620 327134 561240 327218
rect 560620 326898 560652 327134
rect 560888 326898 560972 327134
rect 561208 326898 561240 327134
rect 560620 326866 561240 326898
rect 570260 327454 570880 327486
rect 570260 327218 570292 327454
rect 570528 327218 570612 327454
rect 570848 327218 570880 327454
rect 570260 327134 570880 327218
rect 570260 326898 570292 327134
rect 570528 326898 570612 327134
rect 570848 326898 570880 327134
rect 570260 326866 570880 326898
rect 7844 309454 8464 309486
rect 7844 309218 7876 309454
rect 8112 309218 8196 309454
rect 8432 309218 8464 309454
rect 7844 309134 8464 309218
rect 7844 308898 7876 309134
rect 8112 308898 8196 309134
rect 8432 308898 8464 309134
rect 7844 308866 8464 308898
rect 38000 309454 38620 309486
rect 38000 309218 38032 309454
rect 38268 309218 38352 309454
rect 38588 309218 38620 309454
rect 38000 309134 38620 309218
rect 38000 308898 38032 309134
rect 38268 308898 38352 309134
rect 38588 308898 38620 309134
rect 38000 308866 38620 308898
rect 74000 309454 74620 309486
rect 74000 309218 74032 309454
rect 74268 309218 74352 309454
rect 74588 309218 74620 309454
rect 74000 309134 74620 309218
rect 74000 308898 74032 309134
rect 74268 308898 74352 309134
rect 74588 308898 74620 309134
rect 74000 308866 74620 308898
rect 110000 309454 110620 309486
rect 110000 309218 110032 309454
rect 110268 309218 110352 309454
rect 110588 309218 110620 309454
rect 110000 309134 110620 309218
rect 110000 308898 110032 309134
rect 110268 308898 110352 309134
rect 110588 308898 110620 309134
rect 110000 308866 110620 308898
rect 146000 309454 146620 309486
rect 146000 309218 146032 309454
rect 146268 309218 146352 309454
rect 146588 309218 146620 309454
rect 146000 309134 146620 309218
rect 146000 308898 146032 309134
rect 146268 308898 146352 309134
rect 146588 308898 146620 309134
rect 146000 308866 146620 308898
rect 182000 309454 182620 309486
rect 182000 309218 182032 309454
rect 182268 309218 182352 309454
rect 182588 309218 182620 309454
rect 182000 309134 182620 309218
rect 182000 308898 182032 309134
rect 182268 308898 182352 309134
rect 182588 308898 182620 309134
rect 182000 308866 182620 308898
rect 218000 309454 218620 309486
rect 218000 309218 218032 309454
rect 218268 309218 218352 309454
rect 218588 309218 218620 309454
rect 218000 309134 218620 309218
rect 218000 308898 218032 309134
rect 218268 308898 218352 309134
rect 218588 308898 218620 309134
rect 218000 308866 218620 308898
rect 254000 309454 254620 309486
rect 254000 309218 254032 309454
rect 254268 309218 254352 309454
rect 254588 309218 254620 309454
rect 254000 309134 254620 309218
rect 254000 308898 254032 309134
rect 254268 308898 254352 309134
rect 254588 308898 254620 309134
rect 254000 308866 254620 308898
rect 290000 309454 290620 309486
rect 290000 309218 290032 309454
rect 290268 309218 290352 309454
rect 290588 309218 290620 309454
rect 290000 309134 290620 309218
rect 290000 308898 290032 309134
rect 290268 308898 290352 309134
rect 290588 308898 290620 309134
rect 290000 308866 290620 308898
rect 326000 309454 326620 309486
rect 326000 309218 326032 309454
rect 326268 309218 326352 309454
rect 326588 309218 326620 309454
rect 326000 309134 326620 309218
rect 326000 308898 326032 309134
rect 326268 308898 326352 309134
rect 326588 308898 326620 309134
rect 326000 308866 326620 308898
rect 332293 309454 332653 309486
rect 332293 309218 332355 309454
rect 332591 309218 332653 309454
rect 332293 309134 332653 309218
rect 332293 308898 332355 309134
rect 332591 308898 332653 309134
rect 332293 308866 332653 308898
rect 430769 309454 431129 309486
rect 430769 309218 430831 309454
rect 431067 309218 431129 309454
rect 430769 309134 431129 309218
rect 430769 308898 430831 309134
rect 431067 308898 431129 309134
rect 430769 308866 431129 308898
rect 434000 309454 434620 309486
rect 434000 309218 434032 309454
rect 434268 309218 434352 309454
rect 434588 309218 434620 309454
rect 434000 309134 434620 309218
rect 434000 308898 434032 309134
rect 434268 308898 434352 309134
rect 434588 308898 434620 309134
rect 434000 308866 434620 308898
rect 448249 309454 448609 309486
rect 448249 309218 448311 309454
rect 448547 309218 448609 309454
rect 448249 309134 448609 309218
rect 448249 308898 448311 309134
rect 448547 308898 448609 309134
rect 448249 308866 448609 308898
rect 546725 309454 547085 309486
rect 546725 309218 546787 309454
rect 547023 309218 547085 309454
rect 546725 309134 547085 309218
rect 546725 308898 546787 309134
rect 547023 308898 547085 309134
rect 546725 308866 547085 308898
rect 571500 309454 572120 309486
rect 571500 309218 571532 309454
rect 571768 309218 571852 309454
rect 572088 309218 572120 309454
rect 571500 309134 572120 309218
rect 571500 308898 571532 309134
rect 571768 308898 571852 309134
rect 572088 308898 572120 309134
rect 571500 308866 572120 308898
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect 9084 291454 9704 291486
rect 9084 291218 9116 291454
rect 9352 291218 9436 291454
rect 9672 291218 9704 291454
rect 9084 291134 9704 291218
rect 9084 290898 9116 291134
rect 9352 290898 9436 291134
rect 9672 290898 9704 291134
rect 9084 290866 9704 290898
rect 56620 291454 57240 291486
rect 56620 291218 56652 291454
rect 56888 291218 56972 291454
rect 57208 291218 57240 291454
rect 56620 291134 57240 291218
rect 56620 290898 56652 291134
rect 56888 290898 56972 291134
rect 57208 290898 57240 291134
rect 56620 290866 57240 290898
rect 92620 291454 93240 291486
rect 92620 291218 92652 291454
rect 92888 291218 92972 291454
rect 93208 291218 93240 291454
rect 92620 291134 93240 291218
rect 92620 290898 92652 291134
rect 92888 290898 92972 291134
rect 93208 290898 93240 291134
rect 92620 290866 93240 290898
rect 128620 291454 129240 291486
rect 128620 291218 128652 291454
rect 128888 291218 128972 291454
rect 129208 291218 129240 291454
rect 128620 291134 129240 291218
rect 128620 290898 128652 291134
rect 128888 290898 128972 291134
rect 129208 290898 129240 291134
rect 128620 290866 129240 290898
rect 164620 291454 165240 291486
rect 164620 291218 164652 291454
rect 164888 291218 164972 291454
rect 165208 291218 165240 291454
rect 164620 291134 165240 291218
rect 164620 290898 164652 291134
rect 164888 290898 164972 291134
rect 165208 290898 165240 291134
rect 164620 290866 165240 290898
rect 200620 291454 201240 291486
rect 200620 291218 200652 291454
rect 200888 291218 200972 291454
rect 201208 291218 201240 291454
rect 200620 291134 201240 291218
rect 200620 290898 200652 291134
rect 200888 290898 200972 291134
rect 201208 290898 201240 291134
rect 200620 290866 201240 290898
rect 236620 291454 237240 291486
rect 236620 291218 236652 291454
rect 236888 291218 236972 291454
rect 237208 291218 237240 291454
rect 236620 291134 237240 291218
rect 236620 290898 236652 291134
rect 236888 290898 236972 291134
rect 237208 290898 237240 291134
rect 236620 290866 237240 290898
rect 272620 291454 273240 291486
rect 272620 291218 272652 291454
rect 272888 291218 272972 291454
rect 273208 291218 273240 291454
rect 272620 291134 273240 291218
rect 272620 290898 272652 291134
rect 272888 290898 272972 291134
rect 273208 290898 273240 291134
rect 272620 290866 273240 290898
rect 308620 291454 309240 291486
rect 308620 291218 308652 291454
rect 308888 291218 308972 291454
rect 309208 291218 309240 291454
rect 308620 291134 309240 291218
rect 308620 290898 308652 291134
rect 308888 290898 308972 291134
rect 309208 290898 309240 291134
rect 308620 290866 309240 290898
rect 344620 291454 345240 291486
rect 344620 291218 344652 291454
rect 344888 291218 344972 291454
rect 345208 291218 345240 291454
rect 344620 291134 345240 291218
rect 344620 290898 344652 291134
rect 344888 290898 344972 291134
rect 345208 290898 345240 291134
rect 344620 290866 345240 290898
rect 380620 291454 381240 291486
rect 380620 291218 380652 291454
rect 380888 291218 380972 291454
rect 381208 291218 381240 291454
rect 380620 291134 381240 291218
rect 380620 290898 380652 291134
rect 380888 290898 380972 291134
rect 381208 290898 381240 291134
rect 380620 290866 381240 290898
rect 416620 291454 417240 291486
rect 416620 291218 416652 291454
rect 416888 291218 416972 291454
rect 417208 291218 417240 291454
rect 416620 291134 417240 291218
rect 416620 290898 416652 291134
rect 416888 290898 416972 291134
rect 417208 290898 417240 291134
rect 416620 290866 417240 290898
rect 452620 291454 453240 291486
rect 452620 291218 452652 291454
rect 452888 291218 452972 291454
rect 453208 291218 453240 291454
rect 452620 291134 453240 291218
rect 452620 290898 452652 291134
rect 452888 290898 452972 291134
rect 453208 290898 453240 291134
rect 452620 290866 453240 290898
rect 488620 291454 489240 291486
rect 488620 291218 488652 291454
rect 488888 291218 488972 291454
rect 489208 291218 489240 291454
rect 488620 291134 489240 291218
rect 488620 290898 488652 291134
rect 488888 290898 488972 291134
rect 489208 290898 489240 291134
rect 488620 290866 489240 290898
rect 524620 291454 525240 291486
rect 524620 291218 524652 291454
rect 524888 291218 524972 291454
rect 525208 291218 525240 291454
rect 524620 291134 525240 291218
rect 524620 290898 524652 291134
rect 524888 290898 524972 291134
rect 525208 290898 525240 291134
rect 524620 290866 525240 290898
rect 560620 291454 561240 291486
rect 560620 291218 560652 291454
rect 560888 291218 560972 291454
rect 561208 291218 561240 291454
rect 560620 291134 561240 291218
rect 560620 290898 560652 291134
rect 560888 290898 560972 291134
rect 561208 290898 561240 291134
rect 560620 290866 561240 290898
rect 570260 291454 570880 291486
rect 570260 291218 570292 291454
rect 570528 291218 570612 291454
rect 570848 291218 570880 291454
rect 570260 291134 570880 291218
rect 570260 290898 570292 291134
rect 570528 290898 570612 291134
rect 570848 290898 570880 291134
rect 570260 290866 570880 290898
rect 7844 273454 8464 273486
rect 7844 273218 7876 273454
rect 8112 273218 8196 273454
rect 8432 273218 8464 273454
rect 7844 273134 8464 273218
rect 7844 272898 7876 273134
rect 8112 272898 8196 273134
rect 8432 272898 8464 273134
rect 7844 272866 8464 272898
rect 38000 273454 38620 273486
rect 38000 273218 38032 273454
rect 38268 273218 38352 273454
rect 38588 273218 38620 273454
rect 38000 273134 38620 273218
rect 38000 272898 38032 273134
rect 38268 272898 38352 273134
rect 38588 272898 38620 273134
rect 38000 272866 38620 272898
rect 74000 273454 74620 273486
rect 74000 273218 74032 273454
rect 74268 273218 74352 273454
rect 74588 273218 74620 273454
rect 74000 273134 74620 273218
rect 74000 272898 74032 273134
rect 74268 272898 74352 273134
rect 74588 272898 74620 273134
rect 74000 272866 74620 272898
rect 110000 273454 110620 273486
rect 110000 273218 110032 273454
rect 110268 273218 110352 273454
rect 110588 273218 110620 273454
rect 110000 273134 110620 273218
rect 110000 272898 110032 273134
rect 110268 272898 110352 273134
rect 110588 272898 110620 273134
rect 110000 272866 110620 272898
rect 146000 273454 146620 273486
rect 146000 273218 146032 273454
rect 146268 273218 146352 273454
rect 146588 273218 146620 273454
rect 146000 273134 146620 273218
rect 146000 272898 146032 273134
rect 146268 272898 146352 273134
rect 146588 272898 146620 273134
rect 146000 272866 146620 272898
rect 182000 273454 182620 273486
rect 182000 273218 182032 273454
rect 182268 273218 182352 273454
rect 182588 273218 182620 273454
rect 182000 273134 182620 273218
rect 182000 272898 182032 273134
rect 182268 272898 182352 273134
rect 182588 272898 182620 273134
rect 182000 272866 182620 272898
rect 218000 273454 218620 273486
rect 218000 273218 218032 273454
rect 218268 273218 218352 273454
rect 218588 273218 218620 273454
rect 218000 273134 218620 273218
rect 218000 272898 218032 273134
rect 218268 272898 218352 273134
rect 218588 272898 218620 273134
rect 218000 272866 218620 272898
rect 254000 273454 254620 273486
rect 254000 273218 254032 273454
rect 254268 273218 254352 273454
rect 254588 273218 254620 273454
rect 254000 273134 254620 273218
rect 254000 272898 254032 273134
rect 254268 272898 254352 273134
rect 254588 272898 254620 273134
rect 254000 272866 254620 272898
rect 290000 273454 290620 273486
rect 290000 273218 290032 273454
rect 290268 273218 290352 273454
rect 290588 273218 290620 273454
rect 290000 273134 290620 273218
rect 290000 272898 290032 273134
rect 290268 272898 290352 273134
rect 290588 272898 290620 273134
rect 290000 272866 290620 272898
rect 326000 273454 326620 273486
rect 326000 273218 326032 273454
rect 326268 273218 326352 273454
rect 326588 273218 326620 273454
rect 326000 273134 326620 273218
rect 326000 272898 326032 273134
rect 326268 272898 326352 273134
rect 326588 272898 326620 273134
rect 326000 272866 326620 272898
rect 362000 273454 362620 273486
rect 362000 273218 362032 273454
rect 362268 273218 362352 273454
rect 362588 273218 362620 273454
rect 362000 273134 362620 273218
rect 362000 272898 362032 273134
rect 362268 272898 362352 273134
rect 362588 272898 362620 273134
rect 362000 272866 362620 272898
rect 398000 273454 398620 273486
rect 398000 273218 398032 273454
rect 398268 273218 398352 273454
rect 398588 273218 398620 273454
rect 398000 273134 398620 273218
rect 398000 272898 398032 273134
rect 398268 272898 398352 273134
rect 398588 272898 398620 273134
rect 398000 272866 398620 272898
rect 434000 273454 434620 273486
rect 434000 273218 434032 273454
rect 434268 273218 434352 273454
rect 434588 273218 434620 273454
rect 434000 273134 434620 273218
rect 434000 272898 434032 273134
rect 434268 272898 434352 273134
rect 434588 272898 434620 273134
rect 434000 272866 434620 272898
rect 470000 273454 470620 273486
rect 470000 273218 470032 273454
rect 470268 273218 470352 273454
rect 470588 273218 470620 273454
rect 470000 273134 470620 273218
rect 470000 272898 470032 273134
rect 470268 272898 470352 273134
rect 470588 272898 470620 273134
rect 470000 272866 470620 272898
rect 506000 273454 506620 273486
rect 506000 273218 506032 273454
rect 506268 273218 506352 273454
rect 506588 273218 506620 273454
rect 506000 273134 506620 273218
rect 506000 272898 506032 273134
rect 506268 272898 506352 273134
rect 506588 272898 506620 273134
rect 506000 272866 506620 272898
rect 542000 273454 542620 273486
rect 542000 273218 542032 273454
rect 542268 273218 542352 273454
rect 542588 273218 542620 273454
rect 542000 273134 542620 273218
rect 542000 272898 542032 273134
rect 542268 272898 542352 273134
rect 542588 272898 542620 273134
rect 542000 272866 542620 272898
rect 571500 273454 572120 273486
rect 571500 273218 571532 273454
rect 571768 273218 571852 273454
rect 572088 273218 572120 273454
rect 571500 273134 572120 273218
rect 571500 272898 571532 273134
rect 571768 272898 571852 273134
rect 572088 272898 572120 273134
rect 571500 272866 572120 272898
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect 9084 255454 9704 255486
rect 9084 255218 9116 255454
rect 9352 255218 9436 255454
rect 9672 255218 9704 255454
rect 9084 255134 9704 255218
rect 9084 254898 9116 255134
rect 9352 254898 9436 255134
rect 9672 254898 9704 255134
rect 9084 254866 9704 254898
rect 56620 255454 57240 255486
rect 56620 255218 56652 255454
rect 56888 255218 56972 255454
rect 57208 255218 57240 255454
rect 56620 255134 57240 255218
rect 56620 254898 56652 255134
rect 56888 254898 56972 255134
rect 57208 254898 57240 255134
rect 56620 254866 57240 254898
rect 92620 255454 93240 255486
rect 92620 255218 92652 255454
rect 92888 255218 92972 255454
rect 93208 255218 93240 255454
rect 92620 255134 93240 255218
rect 92620 254898 92652 255134
rect 92888 254898 92972 255134
rect 93208 254898 93240 255134
rect 92620 254866 93240 254898
rect 128620 255454 129240 255486
rect 128620 255218 128652 255454
rect 128888 255218 128972 255454
rect 129208 255218 129240 255454
rect 128620 255134 129240 255218
rect 128620 254898 128652 255134
rect 128888 254898 128972 255134
rect 129208 254898 129240 255134
rect 128620 254866 129240 254898
rect 164620 255454 165240 255486
rect 164620 255218 164652 255454
rect 164888 255218 164972 255454
rect 165208 255218 165240 255454
rect 164620 255134 165240 255218
rect 164620 254898 164652 255134
rect 164888 254898 164972 255134
rect 165208 254898 165240 255134
rect 164620 254866 165240 254898
rect 200620 255454 201240 255486
rect 200620 255218 200652 255454
rect 200888 255218 200972 255454
rect 201208 255218 201240 255454
rect 200620 255134 201240 255218
rect 200620 254898 200652 255134
rect 200888 254898 200972 255134
rect 201208 254898 201240 255134
rect 200620 254866 201240 254898
rect 236620 255454 237240 255486
rect 236620 255218 236652 255454
rect 236888 255218 236972 255454
rect 237208 255218 237240 255454
rect 236620 255134 237240 255218
rect 236620 254898 236652 255134
rect 236888 254898 236972 255134
rect 237208 254898 237240 255134
rect 236620 254866 237240 254898
rect 272620 255454 273240 255486
rect 272620 255218 272652 255454
rect 272888 255218 272972 255454
rect 273208 255218 273240 255454
rect 272620 255134 273240 255218
rect 272620 254898 272652 255134
rect 272888 254898 272972 255134
rect 273208 254898 273240 255134
rect 272620 254866 273240 254898
rect 308620 255454 309240 255486
rect 308620 255218 308652 255454
rect 308888 255218 308972 255454
rect 309208 255218 309240 255454
rect 308620 255134 309240 255218
rect 308620 254898 308652 255134
rect 308888 254898 308972 255134
rect 309208 254898 309240 255134
rect 308620 254866 309240 254898
rect 344620 255454 345240 255486
rect 344620 255218 344652 255454
rect 344888 255218 344972 255454
rect 345208 255218 345240 255454
rect 344620 255134 345240 255218
rect 344620 254898 344652 255134
rect 344888 254898 344972 255134
rect 345208 254898 345240 255134
rect 344620 254866 345240 254898
rect 380620 255454 381240 255486
rect 380620 255218 380652 255454
rect 380888 255218 380972 255454
rect 381208 255218 381240 255454
rect 380620 255134 381240 255218
rect 380620 254898 380652 255134
rect 380888 254898 380972 255134
rect 381208 254898 381240 255134
rect 380620 254866 381240 254898
rect 416620 255454 417240 255486
rect 416620 255218 416652 255454
rect 416888 255218 416972 255454
rect 417208 255218 417240 255454
rect 416620 255134 417240 255218
rect 416620 254898 416652 255134
rect 416888 254898 416972 255134
rect 417208 254898 417240 255134
rect 416620 254866 417240 254898
rect 452620 255454 453240 255486
rect 452620 255218 452652 255454
rect 452888 255218 452972 255454
rect 453208 255218 453240 255454
rect 452620 255134 453240 255218
rect 452620 254898 452652 255134
rect 452888 254898 452972 255134
rect 453208 254898 453240 255134
rect 452620 254866 453240 254898
rect 488620 255454 489240 255486
rect 488620 255218 488652 255454
rect 488888 255218 488972 255454
rect 489208 255218 489240 255454
rect 488620 255134 489240 255218
rect 488620 254898 488652 255134
rect 488888 254898 488972 255134
rect 489208 254898 489240 255134
rect 488620 254866 489240 254898
rect 524620 255454 525240 255486
rect 524620 255218 524652 255454
rect 524888 255218 524972 255454
rect 525208 255218 525240 255454
rect 524620 255134 525240 255218
rect 524620 254898 524652 255134
rect 524888 254898 524972 255134
rect 525208 254898 525240 255134
rect 524620 254866 525240 254898
rect 560620 255454 561240 255486
rect 560620 255218 560652 255454
rect 560888 255218 560972 255454
rect 561208 255218 561240 255454
rect 560620 255134 561240 255218
rect 560620 254898 560652 255134
rect 560888 254898 560972 255134
rect 561208 254898 561240 255134
rect 560620 254866 561240 254898
rect 570260 255454 570880 255486
rect 570260 255218 570292 255454
rect 570528 255218 570612 255454
rect 570848 255218 570880 255454
rect 570260 255134 570880 255218
rect 570260 254898 570292 255134
rect 570528 254898 570612 255134
rect 570848 254898 570880 255134
rect 570260 254866 570880 254898
rect 7844 237454 8464 237486
rect 7844 237218 7876 237454
rect 8112 237218 8196 237454
rect 8432 237218 8464 237454
rect 7844 237134 8464 237218
rect 7844 236898 7876 237134
rect 8112 236898 8196 237134
rect 8432 236898 8464 237134
rect 7844 236866 8464 236898
rect 38000 237454 38620 237486
rect 38000 237218 38032 237454
rect 38268 237218 38352 237454
rect 38588 237218 38620 237454
rect 38000 237134 38620 237218
rect 38000 236898 38032 237134
rect 38268 236898 38352 237134
rect 38588 236898 38620 237134
rect 38000 236866 38620 236898
rect 74000 237454 74620 237486
rect 74000 237218 74032 237454
rect 74268 237218 74352 237454
rect 74588 237218 74620 237454
rect 74000 237134 74620 237218
rect 74000 236898 74032 237134
rect 74268 236898 74352 237134
rect 74588 236898 74620 237134
rect 74000 236866 74620 236898
rect 110000 237454 110620 237486
rect 110000 237218 110032 237454
rect 110268 237218 110352 237454
rect 110588 237218 110620 237454
rect 110000 237134 110620 237218
rect 110000 236898 110032 237134
rect 110268 236898 110352 237134
rect 110588 236898 110620 237134
rect 110000 236866 110620 236898
rect 146000 237454 146620 237486
rect 146000 237218 146032 237454
rect 146268 237218 146352 237454
rect 146588 237218 146620 237454
rect 146000 237134 146620 237218
rect 146000 236898 146032 237134
rect 146268 236898 146352 237134
rect 146588 236898 146620 237134
rect 146000 236866 146620 236898
rect 182000 237454 182620 237486
rect 182000 237218 182032 237454
rect 182268 237218 182352 237454
rect 182588 237218 182620 237454
rect 182000 237134 182620 237218
rect 182000 236898 182032 237134
rect 182268 236898 182352 237134
rect 182588 236898 182620 237134
rect 182000 236866 182620 236898
rect 218000 237454 218620 237486
rect 218000 237218 218032 237454
rect 218268 237218 218352 237454
rect 218588 237218 218620 237454
rect 218000 237134 218620 237218
rect 218000 236898 218032 237134
rect 218268 236898 218352 237134
rect 218588 236898 218620 237134
rect 218000 236866 218620 236898
rect 254000 237454 254620 237486
rect 254000 237218 254032 237454
rect 254268 237218 254352 237454
rect 254588 237218 254620 237454
rect 254000 237134 254620 237218
rect 254000 236898 254032 237134
rect 254268 236898 254352 237134
rect 254588 236898 254620 237134
rect 254000 236866 254620 236898
rect 290000 237454 290620 237486
rect 290000 237218 290032 237454
rect 290268 237218 290352 237454
rect 290588 237218 290620 237454
rect 290000 237134 290620 237218
rect 290000 236898 290032 237134
rect 290268 236898 290352 237134
rect 290588 236898 290620 237134
rect 290000 236866 290620 236898
rect 326000 237454 326620 237486
rect 326000 237218 326032 237454
rect 326268 237218 326352 237454
rect 326588 237218 326620 237454
rect 326000 237134 326620 237218
rect 326000 236898 326032 237134
rect 326268 236898 326352 237134
rect 326588 236898 326620 237134
rect 326000 236866 326620 236898
rect 362000 237454 362620 237486
rect 362000 237218 362032 237454
rect 362268 237218 362352 237454
rect 362588 237218 362620 237454
rect 362000 237134 362620 237218
rect 362000 236898 362032 237134
rect 362268 236898 362352 237134
rect 362588 236898 362620 237134
rect 362000 236866 362620 236898
rect 398000 237454 398620 237486
rect 398000 237218 398032 237454
rect 398268 237218 398352 237454
rect 398588 237218 398620 237454
rect 398000 237134 398620 237218
rect 398000 236898 398032 237134
rect 398268 236898 398352 237134
rect 398588 236898 398620 237134
rect 398000 236866 398620 236898
rect 434000 237454 434620 237486
rect 434000 237218 434032 237454
rect 434268 237218 434352 237454
rect 434588 237218 434620 237454
rect 434000 237134 434620 237218
rect 434000 236898 434032 237134
rect 434268 236898 434352 237134
rect 434588 236898 434620 237134
rect 434000 236866 434620 236898
rect 470000 237454 470620 237486
rect 470000 237218 470032 237454
rect 470268 237218 470352 237454
rect 470588 237218 470620 237454
rect 470000 237134 470620 237218
rect 470000 236898 470032 237134
rect 470268 236898 470352 237134
rect 470588 236898 470620 237134
rect 470000 236866 470620 236898
rect 506000 237454 506620 237486
rect 506000 237218 506032 237454
rect 506268 237218 506352 237454
rect 506588 237218 506620 237454
rect 506000 237134 506620 237218
rect 506000 236898 506032 237134
rect 506268 236898 506352 237134
rect 506588 236898 506620 237134
rect 506000 236866 506620 236898
rect 542000 237454 542620 237486
rect 542000 237218 542032 237454
rect 542268 237218 542352 237454
rect 542588 237218 542620 237454
rect 542000 237134 542620 237218
rect 542000 236898 542032 237134
rect 542268 236898 542352 237134
rect 542588 236898 542620 237134
rect 542000 236866 542620 236898
rect 571500 237454 572120 237486
rect 571500 237218 571532 237454
rect 571768 237218 571852 237454
rect 572088 237218 572120 237454
rect 571500 237134 572120 237218
rect 571500 236898 571532 237134
rect 571768 236898 571852 237134
rect 572088 236898 572120 237134
rect 571500 236866 572120 236898
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect 9084 219454 9704 219486
rect 9084 219218 9116 219454
rect 9352 219218 9436 219454
rect 9672 219218 9704 219454
rect 9084 219134 9704 219218
rect 9084 218898 9116 219134
rect 9352 218898 9436 219134
rect 9672 218898 9704 219134
rect 9084 218866 9704 218898
rect 56620 219454 57240 219486
rect 56620 219218 56652 219454
rect 56888 219218 56972 219454
rect 57208 219218 57240 219454
rect 56620 219134 57240 219218
rect 56620 218898 56652 219134
rect 56888 218898 56972 219134
rect 57208 218898 57240 219134
rect 56620 218866 57240 218898
rect 92620 219454 93240 219486
rect 92620 219218 92652 219454
rect 92888 219218 92972 219454
rect 93208 219218 93240 219454
rect 92620 219134 93240 219218
rect 92620 218898 92652 219134
rect 92888 218898 92972 219134
rect 93208 218898 93240 219134
rect 92620 218866 93240 218898
rect 128620 219454 129240 219486
rect 128620 219218 128652 219454
rect 128888 219218 128972 219454
rect 129208 219218 129240 219454
rect 128620 219134 129240 219218
rect 128620 218898 128652 219134
rect 128888 218898 128972 219134
rect 129208 218898 129240 219134
rect 128620 218866 129240 218898
rect 164620 219454 165240 219486
rect 164620 219218 164652 219454
rect 164888 219218 164972 219454
rect 165208 219218 165240 219454
rect 164620 219134 165240 219218
rect 164620 218898 164652 219134
rect 164888 218898 164972 219134
rect 165208 218898 165240 219134
rect 164620 218866 165240 218898
rect 200620 219454 201240 219486
rect 200620 219218 200652 219454
rect 200888 219218 200972 219454
rect 201208 219218 201240 219454
rect 200620 219134 201240 219218
rect 200620 218898 200652 219134
rect 200888 218898 200972 219134
rect 201208 218898 201240 219134
rect 200620 218866 201240 218898
rect 236620 219454 237240 219486
rect 236620 219218 236652 219454
rect 236888 219218 236972 219454
rect 237208 219218 237240 219454
rect 236620 219134 237240 219218
rect 236620 218898 236652 219134
rect 236888 218898 236972 219134
rect 237208 218898 237240 219134
rect 236620 218866 237240 218898
rect 272620 219454 273240 219486
rect 272620 219218 272652 219454
rect 272888 219218 272972 219454
rect 273208 219218 273240 219454
rect 272620 219134 273240 219218
rect 272620 218898 272652 219134
rect 272888 218898 272972 219134
rect 273208 218898 273240 219134
rect 272620 218866 273240 218898
rect 308620 219454 309240 219486
rect 308620 219218 308652 219454
rect 308888 219218 308972 219454
rect 309208 219218 309240 219454
rect 308620 219134 309240 219218
rect 308620 218898 308652 219134
rect 308888 218898 308972 219134
rect 309208 218898 309240 219134
rect 308620 218866 309240 218898
rect 344620 219454 345240 219486
rect 344620 219218 344652 219454
rect 344888 219218 344972 219454
rect 345208 219218 345240 219454
rect 344620 219134 345240 219218
rect 344620 218898 344652 219134
rect 344888 218898 344972 219134
rect 345208 218898 345240 219134
rect 344620 218866 345240 218898
rect 380620 219454 381240 219486
rect 380620 219218 380652 219454
rect 380888 219218 380972 219454
rect 381208 219218 381240 219454
rect 380620 219134 381240 219218
rect 380620 218898 380652 219134
rect 380888 218898 380972 219134
rect 381208 218898 381240 219134
rect 380620 218866 381240 218898
rect 416620 219454 417240 219486
rect 416620 219218 416652 219454
rect 416888 219218 416972 219454
rect 417208 219218 417240 219454
rect 416620 219134 417240 219218
rect 416620 218898 416652 219134
rect 416888 218898 416972 219134
rect 417208 218898 417240 219134
rect 416620 218866 417240 218898
rect 452620 219454 453240 219486
rect 452620 219218 452652 219454
rect 452888 219218 452972 219454
rect 453208 219218 453240 219454
rect 452620 219134 453240 219218
rect 452620 218898 452652 219134
rect 452888 218898 452972 219134
rect 453208 218898 453240 219134
rect 452620 218866 453240 218898
rect 488620 219454 489240 219486
rect 488620 219218 488652 219454
rect 488888 219218 488972 219454
rect 489208 219218 489240 219454
rect 488620 219134 489240 219218
rect 488620 218898 488652 219134
rect 488888 218898 488972 219134
rect 489208 218898 489240 219134
rect 488620 218866 489240 218898
rect 524620 219454 525240 219486
rect 524620 219218 524652 219454
rect 524888 219218 524972 219454
rect 525208 219218 525240 219454
rect 524620 219134 525240 219218
rect 524620 218898 524652 219134
rect 524888 218898 524972 219134
rect 525208 218898 525240 219134
rect 524620 218866 525240 218898
rect 560620 219454 561240 219486
rect 560620 219218 560652 219454
rect 560888 219218 560972 219454
rect 561208 219218 561240 219454
rect 560620 219134 561240 219218
rect 560620 218898 560652 219134
rect 560888 218898 560972 219134
rect 561208 218898 561240 219134
rect 560620 218866 561240 218898
rect 570260 219454 570880 219486
rect 570260 219218 570292 219454
rect 570528 219218 570612 219454
rect 570848 219218 570880 219454
rect 570260 219134 570880 219218
rect 570260 218898 570292 219134
rect 570528 218898 570612 219134
rect 570848 218898 570880 219134
rect 570260 218866 570880 218898
rect 7844 201454 8464 201486
rect 7844 201218 7876 201454
rect 8112 201218 8196 201454
rect 8432 201218 8464 201454
rect 7844 201134 8464 201218
rect 7844 200898 7876 201134
rect 8112 200898 8196 201134
rect 8432 200898 8464 201134
rect 7844 200866 8464 200898
rect 38000 201454 38620 201486
rect 38000 201218 38032 201454
rect 38268 201218 38352 201454
rect 38588 201218 38620 201454
rect 38000 201134 38620 201218
rect 38000 200898 38032 201134
rect 38268 200898 38352 201134
rect 38588 200898 38620 201134
rect 38000 200866 38620 200898
rect 74000 201454 74620 201486
rect 74000 201218 74032 201454
rect 74268 201218 74352 201454
rect 74588 201218 74620 201454
rect 74000 201134 74620 201218
rect 74000 200898 74032 201134
rect 74268 200898 74352 201134
rect 74588 200898 74620 201134
rect 74000 200866 74620 200898
rect 110000 201454 110620 201486
rect 110000 201218 110032 201454
rect 110268 201218 110352 201454
rect 110588 201218 110620 201454
rect 110000 201134 110620 201218
rect 110000 200898 110032 201134
rect 110268 200898 110352 201134
rect 110588 200898 110620 201134
rect 110000 200866 110620 200898
rect 146000 201454 146620 201486
rect 146000 201218 146032 201454
rect 146268 201218 146352 201454
rect 146588 201218 146620 201454
rect 146000 201134 146620 201218
rect 146000 200898 146032 201134
rect 146268 200898 146352 201134
rect 146588 200898 146620 201134
rect 146000 200866 146620 200898
rect 182000 201454 182620 201486
rect 182000 201218 182032 201454
rect 182268 201218 182352 201454
rect 182588 201218 182620 201454
rect 182000 201134 182620 201218
rect 182000 200898 182032 201134
rect 182268 200898 182352 201134
rect 182588 200898 182620 201134
rect 182000 200866 182620 200898
rect 218000 201454 218620 201486
rect 218000 201218 218032 201454
rect 218268 201218 218352 201454
rect 218588 201218 218620 201454
rect 218000 201134 218620 201218
rect 218000 200898 218032 201134
rect 218268 200898 218352 201134
rect 218588 200898 218620 201134
rect 218000 200866 218620 200898
rect 254000 201454 254620 201486
rect 254000 201218 254032 201454
rect 254268 201218 254352 201454
rect 254588 201218 254620 201454
rect 254000 201134 254620 201218
rect 254000 200898 254032 201134
rect 254268 200898 254352 201134
rect 254588 200898 254620 201134
rect 254000 200866 254620 200898
rect 290000 201454 290620 201486
rect 290000 201218 290032 201454
rect 290268 201218 290352 201454
rect 290588 201218 290620 201454
rect 290000 201134 290620 201218
rect 290000 200898 290032 201134
rect 290268 200898 290352 201134
rect 290588 200898 290620 201134
rect 290000 200866 290620 200898
rect 326000 201454 326620 201486
rect 326000 201218 326032 201454
rect 326268 201218 326352 201454
rect 326588 201218 326620 201454
rect 326000 201134 326620 201218
rect 326000 200898 326032 201134
rect 326268 200898 326352 201134
rect 326588 200898 326620 201134
rect 326000 200866 326620 200898
rect 362000 201454 362620 201486
rect 362000 201218 362032 201454
rect 362268 201218 362352 201454
rect 362588 201218 362620 201454
rect 362000 201134 362620 201218
rect 362000 200898 362032 201134
rect 362268 200898 362352 201134
rect 362588 200898 362620 201134
rect 362000 200866 362620 200898
rect 398000 201454 398620 201486
rect 398000 201218 398032 201454
rect 398268 201218 398352 201454
rect 398588 201218 398620 201454
rect 398000 201134 398620 201218
rect 398000 200898 398032 201134
rect 398268 200898 398352 201134
rect 398588 200898 398620 201134
rect 398000 200866 398620 200898
rect 434000 201454 434620 201486
rect 434000 201218 434032 201454
rect 434268 201218 434352 201454
rect 434588 201218 434620 201454
rect 434000 201134 434620 201218
rect 434000 200898 434032 201134
rect 434268 200898 434352 201134
rect 434588 200898 434620 201134
rect 434000 200866 434620 200898
rect 470000 201454 470620 201486
rect 470000 201218 470032 201454
rect 470268 201218 470352 201454
rect 470588 201218 470620 201454
rect 470000 201134 470620 201218
rect 470000 200898 470032 201134
rect 470268 200898 470352 201134
rect 470588 200898 470620 201134
rect 470000 200866 470620 200898
rect 506000 201454 506620 201486
rect 506000 201218 506032 201454
rect 506268 201218 506352 201454
rect 506588 201218 506620 201454
rect 506000 201134 506620 201218
rect 506000 200898 506032 201134
rect 506268 200898 506352 201134
rect 506588 200898 506620 201134
rect 506000 200866 506620 200898
rect 542000 201454 542620 201486
rect 542000 201218 542032 201454
rect 542268 201218 542352 201454
rect 542588 201218 542620 201454
rect 542000 201134 542620 201218
rect 542000 200898 542032 201134
rect 542268 200898 542352 201134
rect 542588 200898 542620 201134
rect 542000 200866 542620 200898
rect 571500 201454 572120 201486
rect 571500 201218 571532 201454
rect 571768 201218 571852 201454
rect 572088 201218 572120 201454
rect 571500 201134 572120 201218
rect 571500 200898 571532 201134
rect 571768 200898 571852 201134
rect 572088 200898 572120 201134
rect 571500 200866 572120 200898
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect 9084 183454 9704 183486
rect 9084 183218 9116 183454
rect 9352 183218 9436 183454
rect 9672 183218 9704 183454
rect 9084 183134 9704 183218
rect 9084 182898 9116 183134
rect 9352 182898 9436 183134
rect 9672 182898 9704 183134
rect 9084 182866 9704 182898
rect 56620 183454 57240 183486
rect 56620 183218 56652 183454
rect 56888 183218 56972 183454
rect 57208 183218 57240 183454
rect 56620 183134 57240 183218
rect 56620 182898 56652 183134
rect 56888 182898 56972 183134
rect 57208 182898 57240 183134
rect 56620 182866 57240 182898
rect 92620 183454 93240 183486
rect 92620 183218 92652 183454
rect 92888 183218 92972 183454
rect 93208 183218 93240 183454
rect 92620 183134 93240 183218
rect 92620 182898 92652 183134
rect 92888 182898 92972 183134
rect 93208 182898 93240 183134
rect 92620 182866 93240 182898
rect 128620 183454 129240 183486
rect 128620 183218 128652 183454
rect 128888 183218 128972 183454
rect 129208 183218 129240 183454
rect 128620 183134 129240 183218
rect 128620 182898 128652 183134
rect 128888 182898 128972 183134
rect 129208 182898 129240 183134
rect 128620 182866 129240 182898
rect 164620 183454 165240 183486
rect 164620 183218 164652 183454
rect 164888 183218 164972 183454
rect 165208 183218 165240 183454
rect 164620 183134 165240 183218
rect 164620 182898 164652 183134
rect 164888 182898 164972 183134
rect 165208 182898 165240 183134
rect 164620 182866 165240 182898
rect 200620 183454 201240 183486
rect 200620 183218 200652 183454
rect 200888 183218 200972 183454
rect 201208 183218 201240 183454
rect 200620 183134 201240 183218
rect 200620 182898 200652 183134
rect 200888 182898 200972 183134
rect 201208 182898 201240 183134
rect 200620 182866 201240 182898
rect 236620 183454 237240 183486
rect 236620 183218 236652 183454
rect 236888 183218 236972 183454
rect 237208 183218 237240 183454
rect 236620 183134 237240 183218
rect 236620 182898 236652 183134
rect 236888 182898 236972 183134
rect 237208 182898 237240 183134
rect 236620 182866 237240 182898
rect 272620 183454 273240 183486
rect 272620 183218 272652 183454
rect 272888 183218 272972 183454
rect 273208 183218 273240 183454
rect 272620 183134 273240 183218
rect 272620 182898 272652 183134
rect 272888 182898 272972 183134
rect 273208 182898 273240 183134
rect 272620 182866 273240 182898
rect 308620 183454 309240 183486
rect 308620 183218 308652 183454
rect 308888 183218 308972 183454
rect 309208 183218 309240 183454
rect 308620 183134 309240 183218
rect 308620 182898 308652 183134
rect 308888 182898 308972 183134
rect 309208 182898 309240 183134
rect 308620 182866 309240 182898
rect 344620 183454 345240 183486
rect 344620 183218 344652 183454
rect 344888 183218 344972 183454
rect 345208 183218 345240 183454
rect 344620 183134 345240 183218
rect 344620 182898 344652 183134
rect 344888 182898 344972 183134
rect 345208 182898 345240 183134
rect 344620 182866 345240 182898
rect 380620 183454 381240 183486
rect 380620 183218 380652 183454
rect 380888 183218 380972 183454
rect 381208 183218 381240 183454
rect 380620 183134 381240 183218
rect 380620 182898 380652 183134
rect 380888 182898 380972 183134
rect 381208 182898 381240 183134
rect 380620 182866 381240 182898
rect 416620 183454 417240 183486
rect 416620 183218 416652 183454
rect 416888 183218 416972 183454
rect 417208 183218 417240 183454
rect 416620 183134 417240 183218
rect 416620 182898 416652 183134
rect 416888 182898 416972 183134
rect 417208 182898 417240 183134
rect 416620 182866 417240 182898
rect 452620 183454 453240 183486
rect 452620 183218 452652 183454
rect 452888 183218 452972 183454
rect 453208 183218 453240 183454
rect 452620 183134 453240 183218
rect 452620 182898 452652 183134
rect 452888 182898 452972 183134
rect 453208 182898 453240 183134
rect 452620 182866 453240 182898
rect 488620 183454 489240 183486
rect 488620 183218 488652 183454
rect 488888 183218 488972 183454
rect 489208 183218 489240 183454
rect 488620 183134 489240 183218
rect 488620 182898 488652 183134
rect 488888 182898 488972 183134
rect 489208 182898 489240 183134
rect 488620 182866 489240 182898
rect 524620 183454 525240 183486
rect 524620 183218 524652 183454
rect 524888 183218 524972 183454
rect 525208 183218 525240 183454
rect 524620 183134 525240 183218
rect 524620 182898 524652 183134
rect 524888 182898 524972 183134
rect 525208 182898 525240 183134
rect 524620 182866 525240 182898
rect 560620 183454 561240 183486
rect 560620 183218 560652 183454
rect 560888 183218 560972 183454
rect 561208 183218 561240 183454
rect 560620 183134 561240 183218
rect 560620 182898 560652 183134
rect 560888 182898 560972 183134
rect 561208 182898 561240 183134
rect 560620 182866 561240 182898
rect 570260 183454 570880 183486
rect 570260 183218 570292 183454
rect 570528 183218 570612 183454
rect 570848 183218 570880 183454
rect 570260 183134 570880 183218
rect 570260 182898 570292 183134
rect 570528 182898 570612 183134
rect 570848 182898 570880 183134
rect 570260 182866 570880 182898
rect 7844 165454 8464 165486
rect 7844 165218 7876 165454
rect 8112 165218 8196 165454
rect 8432 165218 8464 165454
rect 7844 165134 8464 165218
rect 7844 164898 7876 165134
rect 8112 164898 8196 165134
rect 8432 164898 8464 165134
rect 7844 164866 8464 164898
rect 38000 165454 38620 165486
rect 38000 165218 38032 165454
rect 38268 165218 38352 165454
rect 38588 165218 38620 165454
rect 38000 165134 38620 165218
rect 38000 164898 38032 165134
rect 38268 164898 38352 165134
rect 38588 164898 38620 165134
rect 38000 164866 38620 164898
rect 74000 165454 74620 165486
rect 74000 165218 74032 165454
rect 74268 165218 74352 165454
rect 74588 165218 74620 165454
rect 74000 165134 74620 165218
rect 74000 164898 74032 165134
rect 74268 164898 74352 165134
rect 74588 164898 74620 165134
rect 74000 164866 74620 164898
rect 110000 165454 110620 165486
rect 110000 165218 110032 165454
rect 110268 165218 110352 165454
rect 110588 165218 110620 165454
rect 110000 165134 110620 165218
rect 110000 164898 110032 165134
rect 110268 164898 110352 165134
rect 110588 164898 110620 165134
rect 110000 164866 110620 164898
rect 146000 165454 146620 165486
rect 146000 165218 146032 165454
rect 146268 165218 146352 165454
rect 146588 165218 146620 165454
rect 146000 165134 146620 165218
rect 146000 164898 146032 165134
rect 146268 164898 146352 165134
rect 146588 164898 146620 165134
rect 146000 164866 146620 164898
rect 182000 165454 182620 165486
rect 182000 165218 182032 165454
rect 182268 165218 182352 165454
rect 182588 165218 182620 165454
rect 182000 165134 182620 165218
rect 182000 164898 182032 165134
rect 182268 164898 182352 165134
rect 182588 164898 182620 165134
rect 182000 164866 182620 164898
rect 218000 165454 218620 165486
rect 218000 165218 218032 165454
rect 218268 165218 218352 165454
rect 218588 165218 218620 165454
rect 218000 165134 218620 165218
rect 218000 164898 218032 165134
rect 218268 164898 218352 165134
rect 218588 164898 218620 165134
rect 218000 164866 218620 164898
rect 254000 165454 254620 165486
rect 254000 165218 254032 165454
rect 254268 165218 254352 165454
rect 254588 165218 254620 165454
rect 254000 165134 254620 165218
rect 254000 164898 254032 165134
rect 254268 164898 254352 165134
rect 254588 164898 254620 165134
rect 254000 164866 254620 164898
rect 290000 165454 290620 165486
rect 290000 165218 290032 165454
rect 290268 165218 290352 165454
rect 290588 165218 290620 165454
rect 290000 165134 290620 165218
rect 290000 164898 290032 165134
rect 290268 164898 290352 165134
rect 290588 164898 290620 165134
rect 290000 164866 290620 164898
rect 326000 165454 326620 165486
rect 326000 165218 326032 165454
rect 326268 165218 326352 165454
rect 326588 165218 326620 165454
rect 326000 165134 326620 165218
rect 326000 164898 326032 165134
rect 326268 164898 326352 165134
rect 326588 164898 326620 165134
rect 326000 164866 326620 164898
rect 362000 165454 362620 165486
rect 362000 165218 362032 165454
rect 362268 165218 362352 165454
rect 362588 165218 362620 165454
rect 362000 165134 362620 165218
rect 362000 164898 362032 165134
rect 362268 164898 362352 165134
rect 362588 164898 362620 165134
rect 362000 164866 362620 164898
rect 398000 165454 398620 165486
rect 398000 165218 398032 165454
rect 398268 165218 398352 165454
rect 398588 165218 398620 165454
rect 398000 165134 398620 165218
rect 398000 164898 398032 165134
rect 398268 164898 398352 165134
rect 398588 164898 398620 165134
rect 398000 164866 398620 164898
rect 434000 165454 434620 165486
rect 434000 165218 434032 165454
rect 434268 165218 434352 165454
rect 434588 165218 434620 165454
rect 434000 165134 434620 165218
rect 434000 164898 434032 165134
rect 434268 164898 434352 165134
rect 434588 164898 434620 165134
rect 434000 164866 434620 164898
rect 470000 165454 470620 165486
rect 470000 165218 470032 165454
rect 470268 165218 470352 165454
rect 470588 165218 470620 165454
rect 470000 165134 470620 165218
rect 470000 164898 470032 165134
rect 470268 164898 470352 165134
rect 470588 164898 470620 165134
rect 470000 164866 470620 164898
rect 506000 165454 506620 165486
rect 506000 165218 506032 165454
rect 506268 165218 506352 165454
rect 506588 165218 506620 165454
rect 506000 165134 506620 165218
rect 506000 164898 506032 165134
rect 506268 164898 506352 165134
rect 506588 164898 506620 165134
rect 506000 164866 506620 164898
rect 542000 165454 542620 165486
rect 542000 165218 542032 165454
rect 542268 165218 542352 165454
rect 542588 165218 542620 165454
rect 542000 165134 542620 165218
rect 542000 164898 542032 165134
rect 542268 164898 542352 165134
rect 542588 164898 542620 165134
rect 542000 164866 542620 164898
rect 571500 165454 572120 165486
rect 571500 165218 571532 165454
rect 571768 165218 571852 165454
rect 572088 165218 572120 165454
rect 571500 165134 572120 165218
rect 571500 164898 571532 165134
rect 571768 164898 571852 165134
rect 572088 164898 572120 165134
rect 571500 164866 572120 164898
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect 9084 147454 9704 147486
rect 9084 147218 9116 147454
rect 9352 147218 9436 147454
rect 9672 147218 9704 147454
rect 9084 147134 9704 147218
rect 9084 146898 9116 147134
rect 9352 146898 9436 147134
rect 9672 146898 9704 147134
rect 9084 146866 9704 146898
rect 56620 147454 57240 147486
rect 56620 147218 56652 147454
rect 56888 147218 56972 147454
rect 57208 147218 57240 147454
rect 56620 147134 57240 147218
rect 56620 146898 56652 147134
rect 56888 146898 56972 147134
rect 57208 146898 57240 147134
rect 56620 146866 57240 146898
rect 92620 147454 93240 147486
rect 92620 147218 92652 147454
rect 92888 147218 92972 147454
rect 93208 147218 93240 147454
rect 92620 147134 93240 147218
rect 92620 146898 92652 147134
rect 92888 146898 92972 147134
rect 93208 146898 93240 147134
rect 92620 146866 93240 146898
rect 128620 147454 129240 147486
rect 128620 147218 128652 147454
rect 128888 147218 128972 147454
rect 129208 147218 129240 147454
rect 128620 147134 129240 147218
rect 128620 146898 128652 147134
rect 128888 146898 128972 147134
rect 129208 146898 129240 147134
rect 128620 146866 129240 146898
rect 164620 147454 165240 147486
rect 164620 147218 164652 147454
rect 164888 147218 164972 147454
rect 165208 147218 165240 147454
rect 164620 147134 165240 147218
rect 164620 146898 164652 147134
rect 164888 146898 164972 147134
rect 165208 146898 165240 147134
rect 164620 146866 165240 146898
rect 200620 147454 201240 147486
rect 200620 147218 200652 147454
rect 200888 147218 200972 147454
rect 201208 147218 201240 147454
rect 200620 147134 201240 147218
rect 200620 146898 200652 147134
rect 200888 146898 200972 147134
rect 201208 146898 201240 147134
rect 200620 146866 201240 146898
rect 236620 147454 237240 147486
rect 236620 147218 236652 147454
rect 236888 147218 236972 147454
rect 237208 147218 237240 147454
rect 236620 147134 237240 147218
rect 236620 146898 236652 147134
rect 236888 146898 236972 147134
rect 237208 146898 237240 147134
rect 236620 146866 237240 146898
rect 272620 147454 273240 147486
rect 272620 147218 272652 147454
rect 272888 147218 272972 147454
rect 273208 147218 273240 147454
rect 272620 147134 273240 147218
rect 272620 146898 272652 147134
rect 272888 146898 272972 147134
rect 273208 146898 273240 147134
rect 272620 146866 273240 146898
rect 308620 147454 309240 147486
rect 308620 147218 308652 147454
rect 308888 147218 308972 147454
rect 309208 147218 309240 147454
rect 308620 147134 309240 147218
rect 308620 146898 308652 147134
rect 308888 146898 308972 147134
rect 309208 146898 309240 147134
rect 308620 146866 309240 146898
rect 344620 147454 345240 147486
rect 344620 147218 344652 147454
rect 344888 147218 344972 147454
rect 345208 147218 345240 147454
rect 344620 147134 345240 147218
rect 344620 146898 344652 147134
rect 344888 146898 344972 147134
rect 345208 146898 345240 147134
rect 344620 146866 345240 146898
rect 380620 147454 381240 147486
rect 380620 147218 380652 147454
rect 380888 147218 380972 147454
rect 381208 147218 381240 147454
rect 380620 147134 381240 147218
rect 380620 146898 380652 147134
rect 380888 146898 380972 147134
rect 381208 146898 381240 147134
rect 380620 146866 381240 146898
rect 416620 147454 417240 147486
rect 416620 147218 416652 147454
rect 416888 147218 416972 147454
rect 417208 147218 417240 147454
rect 416620 147134 417240 147218
rect 416620 146898 416652 147134
rect 416888 146898 416972 147134
rect 417208 146898 417240 147134
rect 416620 146866 417240 146898
rect 452620 147454 453240 147486
rect 452620 147218 452652 147454
rect 452888 147218 452972 147454
rect 453208 147218 453240 147454
rect 452620 147134 453240 147218
rect 452620 146898 452652 147134
rect 452888 146898 452972 147134
rect 453208 146898 453240 147134
rect 452620 146866 453240 146898
rect 488620 147454 489240 147486
rect 488620 147218 488652 147454
rect 488888 147218 488972 147454
rect 489208 147218 489240 147454
rect 488620 147134 489240 147218
rect 488620 146898 488652 147134
rect 488888 146898 488972 147134
rect 489208 146898 489240 147134
rect 488620 146866 489240 146898
rect 524620 147454 525240 147486
rect 524620 147218 524652 147454
rect 524888 147218 524972 147454
rect 525208 147218 525240 147454
rect 524620 147134 525240 147218
rect 524620 146898 524652 147134
rect 524888 146898 524972 147134
rect 525208 146898 525240 147134
rect 524620 146866 525240 146898
rect 560620 147454 561240 147486
rect 560620 147218 560652 147454
rect 560888 147218 560972 147454
rect 561208 147218 561240 147454
rect 560620 147134 561240 147218
rect 560620 146898 560652 147134
rect 560888 146898 560972 147134
rect 561208 146898 561240 147134
rect 560620 146866 561240 146898
rect 570260 147454 570880 147486
rect 570260 147218 570292 147454
rect 570528 147218 570612 147454
rect 570848 147218 570880 147454
rect 570260 147134 570880 147218
rect 570260 146898 570292 147134
rect 570528 146898 570612 147134
rect 570848 146898 570880 147134
rect 570260 146866 570880 146898
rect 7844 129454 8464 129486
rect 7844 129218 7876 129454
rect 8112 129218 8196 129454
rect 8432 129218 8464 129454
rect 7844 129134 8464 129218
rect 7844 128898 7876 129134
rect 8112 128898 8196 129134
rect 8432 128898 8464 129134
rect 7844 128866 8464 128898
rect 38000 129454 38620 129486
rect 38000 129218 38032 129454
rect 38268 129218 38352 129454
rect 38588 129218 38620 129454
rect 38000 129134 38620 129218
rect 38000 128898 38032 129134
rect 38268 128898 38352 129134
rect 38588 128898 38620 129134
rect 38000 128866 38620 128898
rect 74000 129454 74620 129486
rect 74000 129218 74032 129454
rect 74268 129218 74352 129454
rect 74588 129218 74620 129454
rect 74000 129134 74620 129218
rect 74000 128898 74032 129134
rect 74268 128898 74352 129134
rect 74588 128898 74620 129134
rect 74000 128866 74620 128898
rect 110000 129454 110620 129486
rect 110000 129218 110032 129454
rect 110268 129218 110352 129454
rect 110588 129218 110620 129454
rect 110000 129134 110620 129218
rect 110000 128898 110032 129134
rect 110268 128898 110352 129134
rect 110588 128898 110620 129134
rect 110000 128866 110620 128898
rect 146000 129454 146620 129486
rect 146000 129218 146032 129454
rect 146268 129218 146352 129454
rect 146588 129218 146620 129454
rect 146000 129134 146620 129218
rect 146000 128898 146032 129134
rect 146268 128898 146352 129134
rect 146588 128898 146620 129134
rect 146000 128866 146620 128898
rect 182000 129454 182620 129486
rect 182000 129218 182032 129454
rect 182268 129218 182352 129454
rect 182588 129218 182620 129454
rect 182000 129134 182620 129218
rect 182000 128898 182032 129134
rect 182268 128898 182352 129134
rect 182588 128898 182620 129134
rect 182000 128866 182620 128898
rect 218000 129454 218620 129486
rect 218000 129218 218032 129454
rect 218268 129218 218352 129454
rect 218588 129218 218620 129454
rect 218000 129134 218620 129218
rect 218000 128898 218032 129134
rect 218268 128898 218352 129134
rect 218588 128898 218620 129134
rect 218000 128866 218620 128898
rect 254000 129454 254620 129486
rect 254000 129218 254032 129454
rect 254268 129218 254352 129454
rect 254588 129218 254620 129454
rect 254000 129134 254620 129218
rect 254000 128898 254032 129134
rect 254268 128898 254352 129134
rect 254588 128898 254620 129134
rect 254000 128866 254620 128898
rect 290000 129454 290620 129486
rect 290000 129218 290032 129454
rect 290268 129218 290352 129454
rect 290588 129218 290620 129454
rect 290000 129134 290620 129218
rect 290000 128898 290032 129134
rect 290268 128898 290352 129134
rect 290588 128898 290620 129134
rect 290000 128866 290620 128898
rect 326000 129454 326620 129486
rect 326000 129218 326032 129454
rect 326268 129218 326352 129454
rect 326588 129218 326620 129454
rect 326000 129134 326620 129218
rect 326000 128898 326032 129134
rect 326268 128898 326352 129134
rect 326588 128898 326620 129134
rect 326000 128866 326620 128898
rect 362000 129454 362620 129486
rect 362000 129218 362032 129454
rect 362268 129218 362352 129454
rect 362588 129218 362620 129454
rect 362000 129134 362620 129218
rect 362000 128898 362032 129134
rect 362268 128898 362352 129134
rect 362588 128898 362620 129134
rect 362000 128866 362620 128898
rect 398000 129454 398620 129486
rect 398000 129218 398032 129454
rect 398268 129218 398352 129454
rect 398588 129218 398620 129454
rect 398000 129134 398620 129218
rect 398000 128898 398032 129134
rect 398268 128898 398352 129134
rect 398588 128898 398620 129134
rect 398000 128866 398620 128898
rect 434000 129454 434620 129486
rect 434000 129218 434032 129454
rect 434268 129218 434352 129454
rect 434588 129218 434620 129454
rect 434000 129134 434620 129218
rect 434000 128898 434032 129134
rect 434268 128898 434352 129134
rect 434588 128898 434620 129134
rect 434000 128866 434620 128898
rect 470000 129454 470620 129486
rect 470000 129218 470032 129454
rect 470268 129218 470352 129454
rect 470588 129218 470620 129454
rect 470000 129134 470620 129218
rect 470000 128898 470032 129134
rect 470268 128898 470352 129134
rect 470588 128898 470620 129134
rect 470000 128866 470620 128898
rect 506000 129454 506620 129486
rect 506000 129218 506032 129454
rect 506268 129218 506352 129454
rect 506588 129218 506620 129454
rect 506000 129134 506620 129218
rect 506000 128898 506032 129134
rect 506268 128898 506352 129134
rect 506588 128898 506620 129134
rect 506000 128866 506620 128898
rect 542000 129454 542620 129486
rect 542000 129218 542032 129454
rect 542268 129218 542352 129454
rect 542588 129218 542620 129454
rect 542000 129134 542620 129218
rect 542000 128898 542032 129134
rect 542268 128898 542352 129134
rect 542588 128898 542620 129134
rect 542000 128866 542620 128898
rect 571500 129454 572120 129486
rect 571500 129218 571532 129454
rect 571768 129218 571852 129454
rect 572088 129218 572120 129454
rect 571500 129134 572120 129218
rect 571500 128898 571532 129134
rect 571768 128898 571852 129134
rect 572088 128898 572120 129134
rect 571500 128866 572120 128898
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect 9084 111454 9704 111486
rect 9084 111218 9116 111454
rect 9352 111218 9436 111454
rect 9672 111218 9704 111454
rect 9084 111134 9704 111218
rect 9084 110898 9116 111134
rect 9352 110898 9436 111134
rect 9672 110898 9704 111134
rect 9084 110866 9704 110898
rect 56620 111454 57240 111486
rect 56620 111218 56652 111454
rect 56888 111218 56972 111454
rect 57208 111218 57240 111454
rect 56620 111134 57240 111218
rect 56620 110898 56652 111134
rect 56888 110898 56972 111134
rect 57208 110898 57240 111134
rect 56620 110866 57240 110898
rect 92620 111454 93240 111486
rect 92620 111218 92652 111454
rect 92888 111218 92972 111454
rect 93208 111218 93240 111454
rect 92620 111134 93240 111218
rect 92620 110898 92652 111134
rect 92888 110898 92972 111134
rect 93208 110898 93240 111134
rect 92620 110866 93240 110898
rect 128620 111454 129240 111486
rect 128620 111218 128652 111454
rect 128888 111218 128972 111454
rect 129208 111218 129240 111454
rect 128620 111134 129240 111218
rect 128620 110898 128652 111134
rect 128888 110898 128972 111134
rect 129208 110898 129240 111134
rect 128620 110866 129240 110898
rect 164620 111454 165240 111486
rect 164620 111218 164652 111454
rect 164888 111218 164972 111454
rect 165208 111218 165240 111454
rect 164620 111134 165240 111218
rect 164620 110898 164652 111134
rect 164888 110898 164972 111134
rect 165208 110898 165240 111134
rect 164620 110866 165240 110898
rect 200620 111454 201240 111486
rect 200620 111218 200652 111454
rect 200888 111218 200972 111454
rect 201208 111218 201240 111454
rect 200620 111134 201240 111218
rect 200620 110898 200652 111134
rect 200888 110898 200972 111134
rect 201208 110898 201240 111134
rect 200620 110866 201240 110898
rect 236620 111454 237240 111486
rect 236620 111218 236652 111454
rect 236888 111218 236972 111454
rect 237208 111218 237240 111454
rect 236620 111134 237240 111218
rect 236620 110898 236652 111134
rect 236888 110898 236972 111134
rect 237208 110898 237240 111134
rect 236620 110866 237240 110898
rect 272620 111454 273240 111486
rect 272620 111218 272652 111454
rect 272888 111218 272972 111454
rect 273208 111218 273240 111454
rect 272620 111134 273240 111218
rect 272620 110898 272652 111134
rect 272888 110898 272972 111134
rect 273208 110898 273240 111134
rect 272620 110866 273240 110898
rect 308620 111454 309240 111486
rect 308620 111218 308652 111454
rect 308888 111218 308972 111454
rect 309208 111218 309240 111454
rect 308620 111134 309240 111218
rect 308620 110898 308652 111134
rect 308888 110898 308972 111134
rect 309208 110898 309240 111134
rect 308620 110866 309240 110898
rect 344620 111454 345240 111486
rect 344620 111218 344652 111454
rect 344888 111218 344972 111454
rect 345208 111218 345240 111454
rect 344620 111134 345240 111218
rect 344620 110898 344652 111134
rect 344888 110898 344972 111134
rect 345208 110898 345240 111134
rect 344620 110866 345240 110898
rect 380620 111454 381240 111486
rect 380620 111218 380652 111454
rect 380888 111218 380972 111454
rect 381208 111218 381240 111454
rect 380620 111134 381240 111218
rect 380620 110898 380652 111134
rect 380888 110898 380972 111134
rect 381208 110898 381240 111134
rect 380620 110866 381240 110898
rect 416620 111454 417240 111486
rect 416620 111218 416652 111454
rect 416888 111218 416972 111454
rect 417208 111218 417240 111454
rect 416620 111134 417240 111218
rect 416620 110898 416652 111134
rect 416888 110898 416972 111134
rect 417208 110898 417240 111134
rect 416620 110866 417240 110898
rect 452620 111454 453240 111486
rect 452620 111218 452652 111454
rect 452888 111218 452972 111454
rect 453208 111218 453240 111454
rect 452620 111134 453240 111218
rect 452620 110898 452652 111134
rect 452888 110898 452972 111134
rect 453208 110898 453240 111134
rect 452620 110866 453240 110898
rect 488620 111454 489240 111486
rect 488620 111218 488652 111454
rect 488888 111218 488972 111454
rect 489208 111218 489240 111454
rect 488620 111134 489240 111218
rect 488620 110898 488652 111134
rect 488888 110898 488972 111134
rect 489208 110898 489240 111134
rect 488620 110866 489240 110898
rect 524620 111454 525240 111486
rect 524620 111218 524652 111454
rect 524888 111218 524972 111454
rect 525208 111218 525240 111454
rect 524620 111134 525240 111218
rect 524620 110898 524652 111134
rect 524888 110898 524972 111134
rect 525208 110898 525240 111134
rect 524620 110866 525240 110898
rect 560620 111454 561240 111486
rect 560620 111218 560652 111454
rect 560888 111218 560972 111454
rect 561208 111218 561240 111454
rect 560620 111134 561240 111218
rect 560620 110898 560652 111134
rect 560888 110898 560972 111134
rect 561208 110898 561240 111134
rect 560620 110866 561240 110898
rect 570260 111454 570880 111486
rect 570260 111218 570292 111454
rect 570528 111218 570612 111454
rect 570848 111218 570880 111454
rect 570260 111134 570880 111218
rect 570260 110898 570292 111134
rect 570528 110898 570612 111134
rect 570848 110898 570880 111134
rect 570260 110866 570880 110898
rect 7844 93454 8464 93486
rect 7844 93218 7876 93454
rect 8112 93218 8196 93454
rect 8432 93218 8464 93454
rect 7844 93134 8464 93218
rect 7844 92898 7876 93134
rect 8112 92898 8196 93134
rect 8432 92898 8464 93134
rect 7844 92866 8464 92898
rect 38000 93454 38620 93486
rect 38000 93218 38032 93454
rect 38268 93218 38352 93454
rect 38588 93218 38620 93454
rect 38000 93134 38620 93218
rect 38000 92898 38032 93134
rect 38268 92898 38352 93134
rect 38588 92898 38620 93134
rect 38000 92866 38620 92898
rect 74000 93454 74620 93486
rect 74000 93218 74032 93454
rect 74268 93218 74352 93454
rect 74588 93218 74620 93454
rect 74000 93134 74620 93218
rect 74000 92898 74032 93134
rect 74268 92898 74352 93134
rect 74588 92898 74620 93134
rect 74000 92866 74620 92898
rect 110000 93454 110620 93486
rect 110000 93218 110032 93454
rect 110268 93218 110352 93454
rect 110588 93218 110620 93454
rect 110000 93134 110620 93218
rect 110000 92898 110032 93134
rect 110268 92898 110352 93134
rect 110588 92898 110620 93134
rect 110000 92866 110620 92898
rect 146000 93454 146620 93486
rect 146000 93218 146032 93454
rect 146268 93218 146352 93454
rect 146588 93218 146620 93454
rect 146000 93134 146620 93218
rect 146000 92898 146032 93134
rect 146268 92898 146352 93134
rect 146588 92898 146620 93134
rect 146000 92866 146620 92898
rect 182000 93454 182620 93486
rect 182000 93218 182032 93454
rect 182268 93218 182352 93454
rect 182588 93218 182620 93454
rect 182000 93134 182620 93218
rect 182000 92898 182032 93134
rect 182268 92898 182352 93134
rect 182588 92898 182620 93134
rect 182000 92866 182620 92898
rect 218000 93454 218620 93486
rect 218000 93218 218032 93454
rect 218268 93218 218352 93454
rect 218588 93218 218620 93454
rect 218000 93134 218620 93218
rect 218000 92898 218032 93134
rect 218268 92898 218352 93134
rect 218588 92898 218620 93134
rect 218000 92866 218620 92898
rect 254000 93454 254620 93486
rect 254000 93218 254032 93454
rect 254268 93218 254352 93454
rect 254588 93218 254620 93454
rect 254000 93134 254620 93218
rect 254000 92898 254032 93134
rect 254268 92898 254352 93134
rect 254588 92898 254620 93134
rect 254000 92866 254620 92898
rect 290000 93454 290620 93486
rect 290000 93218 290032 93454
rect 290268 93218 290352 93454
rect 290588 93218 290620 93454
rect 290000 93134 290620 93218
rect 290000 92898 290032 93134
rect 290268 92898 290352 93134
rect 290588 92898 290620 93134
rect 290000 92866 290620 92898
rect 326000 93454 326620 93486
rect 326000 93218 326032 93454
rect 326268 93218 326352 93454
rect 326588 93218 326620 93454
rect 326000 93134 326620 93218
rect 326000 92898 326032 93134
rect 326268 92898 326352 93134
rect 326588 92898 326620 93134
rect 326000 92866 326620 92898
rect 362000 93454 362620 93486
rect 362000 93218 362032 93454
rect 362268 93218 362352 93454
rect 362588 93218 362620 93454
rect 362000 93134 362620 93218
rect 362000 92898 362032 93134
rect 362268 92898 362352 93134
rect 362588 92898 362620 93134
rect 362000 92866 362620 92898
rect 398000 93454 398620 93486
rect 398000 93218 398032 93454
rect 398268 93218 398352 93454
rect 398588 93218 398620 93454
rect 398000 93134 398620 93218
rect 398000 92898 398032 93134
rect 398268 92898 398352 93134
rect 398588 92898 398620 93134
rect 398000 92866 398620 92898
rect 434000 93454 434620 93486
rect 434000 93218 434032 93454
rect 434268 93218 434352 93454
rect 434588 93218 434620 93454
rect 434000 93134 434620 93218
rect 434000 92898 434032 93134
rect 434268 92898 434352 93134
rect 434588 92898 434620 93134
rect 434000 92866 434620 92898
rect 470000 93454 470620 93486
rect 470000 93218 470032 93454
rect 470268 93218 470352 93454
rect 470588 93218 470620 93454
rect 470000 93134 470620 93218
rect 470000 92898 470032 93134
rect 470268 92898 470352 93134
rect 470588 92898 470620 93134
rect 470000 92866 470620 92898
rect 506000 93454 506620 93486
rect 506000 93218 506032 93454
rect 506268 93218 506352 93454
rect 506588 93218 506620 93454
rect 506000 93134 506620 93218
rect 506000 92898 506032 93134
rect 506268 92898 506352 93134
rect 506588 92898 506620 93134
rect 506000 92866 506620 92898
rect 542000 93454 542620 93486
rect 542000 93218 542032 93454
rect 542268 93218 542352 93454
rect 542588 93218 542620 93454
rect 542000 93134 542620 93218
rect 542000 92898 542032 93134
rect 542268 92898 542352 93134
rect 542588 92898 542620 93134
rect 542000 92866 542620 92898
rect 571500 93454 572120 93486
rect 571500 93218 571532 93454
rect 571768 93218 571852 93454
rect 572088 93218 572120 93454
rect 571500 93134 572120 93218
rect 571500 92898 571532 93134
rect 571768 92898 571852 93134
rect 572088 92898 572120 93134
rect 571500 92866 572120 92898
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect 9084 75454 9704 75486
rect 9084 75218 9116 75454
rect 9352 75218 9436 75454
rect 9672 75218 9704 75454
rect 9084 75134 9704 75218
rect 9084 74898 9116 75134
rect 9352 74898 9436 75134
rect 9672 74898 9704 75134
rect 9084 74866 9704 74898
rect 56620 75454 57240 75486
rect 56620 75218 56652 75454
rect 56888 75218 56972 75454
rect 57208 75218 57240 75454
rect 56620 75134 57240 75218
rect 56620 74898 56652 75134
rect 56888 74898 56972 75134
rect 57208 74898 57240 75134
rect 56620 74866 57240 74898
rect 92620 75454 93240 75486
rect 92620 75218 92652 75454
rect 92888 75218 92972 75454
rect 93208 75218 93240 75454
rect 92620 75134 93240 75218
rect 92620 74898 92652 75134
rect 92888 74898 92972 75134
rect 93208 74898 93240 75134
rect 92620 74866 93240 74898
rect 128620 75454 129240 75486
rect 128620 75218 128652 75454
rect 128888 75218 128972 75454
rect 129208 75218 129240 75454
rect 128620 75134 129240 75218
rect 128620 74898 128652 75134
rect 128888 74898 128972 75134
rect 129208 74898 129240 75134
rect 128620 74866 129240 74898
rect 164620 75454 165240 75486
rect 164620 75218 164652 75454
rect 164888 75218 164972 75454
rect 165208 75218 165240 75454
rect 164620 75134 165240 75218
rect 164620 74898 164652 75134
rect 164888 74898 164972 75134
rect 165208 74898 165240 75134
rect 164620 74866 165240 74898
rect 200620 75454 201240 75486
rect 200620 75218 200652 75454
rect 200888 75218 200972 75454
rect 201208 75218 201240 75454
rect 200620 75134 201240 75218
rect 200620 74898 200652 75134
rect 200888 74898 200972 75134
rect 201208 74898 201240 75134
rect 200620 74866 201240 74898
rect 236620 75454 237240 75486
rect 236620 75218 236652 75454
rect 236888 75218 236972 75454
rect 237208 75218 237240 75454
rect 236620 75134 237240 75218
rect 236620 74898 236652 75134
rect 236888 74898 236972 75134
rect 237208 74898 237240 75134
rect 236620 74866 237240 74898
rect 272620 75454 273240 75486
rect 272620 75218 272652 75454
rect 272888 75218 272972 75454
rect 273208 75218 273240 75454
rect 272620 75134 273240 75218
rect 272620 74898 272652 75134
rect 272888 74898 272972 75134
rect 273208 74898 273240 75134
rect 272620 74866 273240 74898
rect 308620 75454 309240 75486
rect 308620 75218 308652 75454
rect 308888 75218 308972 75454
rect 309208 75218 309240 75454
rect 308620 75134 309240 75218
rect 308620 74898 308652 75134
rect 308888 74898 308972 75134
rect 309208 74898 309240 75134
rect 308620 74866 309240 74898
rect 344620 75454 345240 75486
rect 344620 75218 344652 75454
rect 344888 75218 344972 75454
rect 345208 75218 345240 75454
rect 344620 75134 345240 75218
rect 344620 74898 344652 75134
rect 344888 74898 344972 75134
rect 345208 74898 345240 75134
rect 344620 74866 345240 74898
rect 380620 75454 381240 75486
rect 380620 75218 380652 75454
rect 380888 75218 380972 75454
rect 381208 75218 381240 75454
rect 380620 75134 381240 75218
rect 380620 74898 380652 75134
rect 380888 74898 380972 75134
rect 381208 74898 381240 75134
rect 380620 74866 381240 74898
rect 416620 75454 417240 75486
rect 416620 75218 416652 75454
rect 416888 75218 416972 75454
rect 417208 75218 417240 75454
rect 416620 75134 417240 75218
rect 416620 74898 416652 75134
rect 416888 74898 416972 75134
rect 417208 74898 417240 75134
rect 416620 74866 417240 74898
rect 452620 75454 453240 75486
rect 452620 75218 452652 75454
rect 452888 75218 452972 75454
rect 453208 75218 453240 75454
rect 452620 75134 453240 75218
rect 452620 74898 452652 75134
rect 452888 74898 452972 75134
rect 453208 74898 453240 75134
rect 452620 74866 453240 74898
rect 488620 75454 489240 75486
rect 488620 75218 488652 75454
rect 488888 75218 488972 75454
rect 489208 75218 489240 75454
rect 488620 75134 489240 75218
rect 488620 74898 488652 75134
rect 488888 74898 488972 75134
rect 489208 74898 489240 75134
rect 488620 74866 489240 74898
rect 524620 75454 525240 75486
rect 524620 75218 524652 75454
rect 524888 75218 524972 75454
rect 525208 75218 525240 75454
rect 524620 75134 525240 75218
rect 524620 74898 524652 75134
rect 524888 74898 524972 75134
rect 525208 74898 525240 75134
rect 524620 74866 525240 74898
rect 560620 75454 561240 75486
rect 560620 75218 560652 75454
rect 560888 75218 560972 75454
rect 561208 75218 561240 75454
rect 560620 75134 561240 75218
rect 560620 74898 560652 75134
rect 560888 74898 560972 75134
rect 561208 74898 561240 75134
rect 560620 74866 561240 74898
rect 570260 75454 570880 75486
rect 570260 75218 570292 75454
rect 570528 75218 570612 75454
rect 570848 75218 570880 75454
rect 570260 75134 570880 75218
rect 570260 74898 570292 75134
rect 570528 74898 570612 75134
rect 570848 74898 570880 75134
rect 570260 74866 570880 74898
rect 7844 57454 8464 57486
rect 7844 57218 7876 57454
rect 8112 57218 8196 57454
rect 8432 57218 8464 57454
rect 7844 57134 8464 57218
rect 7844 56898 7876 57134
rect 8112 56898 8196 57134
rect 8432 56898 8464 57134
rect 7844 56866 8464 56898
rect 38000 57454 38620 57486
rect 38000 57218 38032 57454
rect 38268 57218 38352 57454
rect 38588 57218 38620 57454
rect 38000 57134 38620 57218
rect 38000 56898 38032 57134
rect 38268 56898 38352 57134
rect 38588 56898 38620 57134
rect 38000 56866 38620 56898
rect 74000 57454 74620 57486
rect 74000 57218 74032 57454
rect 74268 57218 74352 57454
rect 74588 57218 74620 57454
rect 74000 57134 74620 57218
rect 74000 56898 74032 57134
rect 74268 56898 74352 57134
rect 74588 56898 74620 57134
rect 74000 56866 74620 56898
rect 110000 57454 110620 57486
rect 110000 57218 110032 57454
rect 110268 57218 110352 57454
rect 110588 57218 110620 57454
rect 110000 57134 110620 57218
rect 110000 56898 110032 57134
rect 110268 56898 110352 57134
rect 110588 56898 110620 57134
rect 110000 56866 110620 56898
rect 146000 57454 146620 57486
rect 146000 57218 146032 57454
rect 146268 57218 146352 57454
rect 146588 57218 146620 57454
rect 146000 57134 146620 57218
rect 146000 56898 146032 57134
rect 146268 56898 146352 57134
rect 146588 56898 146620 57134
rect 146000 56866 146620 56898
rect 182000 57454 182620 57486
rect 182000 57218 182032 57454
rect 182268 57218 182352 57454
rect 182588 57218 182620 57454
rect 182000 57134 182620 57218
rect 182000 56898 182032 57134
rect 182268 56898 182352 57134
rect 182588 56898 182620 57134
rect 182000 56866 182620 56898
rect 218000 57454 218620 57486
rect 218000 57218 218032 57454
rect 218268 57218 218352 57454
rect 218588 57218 218620 57454
rect 218000 57134 218620 57218
rect 218000 56898 218032 57134
rect 218268 56898 218352 57134
rect 218588 56898 218620 57134
rect 218000 56866 218620 56898
rect 254000 57454 254620 57486
rect 254000 57218 254032 57454
rect 254268 57218 254352 57454
rect 254588 57218 254620 57454
rect 254000 57134 254620 57218
rect 254000 56898 254032 57134
rect 254268 56898 254352 57134
rect 254588 56898 254620 57134
rect 254000 56866 254620 56898
rect 290000 57454 290620 57486
rect 290000 57218 290032 57454
rect 290268 57218 290352 57454
rect 290588 57218 290620 57454
rect 290000 57134 290620 57218
rect 290000 56898 290032 57134
rect 290268 56898 290352 57134
rect 290588 56898 290620 57134
rect 290000 56866 290620 56898
rect 326000 57454 326620 57486
rect 326000 57218 326032 57454
rect 326268 57218 326352 57454
rect 326588 57218 326620 57454
rect 326000 57134 326620 57218
rect 326000 56898 326032 57134
rect 326268 56898 326352 57134
rect 326588 56898 326620 57134
rect 326000 56866 326620 56898
rect 362000 57454 362620 57486
rect 362000 57218 362032 57454
rect 362268 57218 362352 57454
rect 362588 57218 362620 57454
rect 362000 57134 362620 57218
rect 362000 56898 362032 57134
rect 362268 56898 362352 57134
rect 362588 56898 362620 57134
rect 362000 56866 362620 56898
rect 398000 57454 398620 57486
rect 398000 57218 398032 57454
rect 398268 57218 398352 57454
rect 398588 57218 398620 57454
rect 398000 57134 398620 57218
rect 398000 56898 398032 57134
rect 398268 56898 398352 57134
rect 398588 56898 398620 57134
rect 398000 56866 398620 56898
rect 434000 57454 434620 57486
rect 434000 57218 434032 57454
rect 434268 57218 434352 57454
rect 434588 57218 434620 57454
rect 434000 57134 434620 57218
rect 434000 56898 434032 57134
rect 434268 56898 434352 57134
rect 434588 56898 434620 57134
rect 434000 56866 434620 56898
rect 470000 57454 470620 57486
rect 470000 57218 470032 57454
rect 470268 57218 470352 57454
rect 470588 57218 470620 57454
rect 470000 57134 470620 57218
rect 470000 56898 470032 57134
rect 470268 56898 470352 57134
rect 470588 56898 470620 57134
rect 470000 56866 470620 56898
rect 506000 57454 506620 57486
rect 506000 57218 506032 57454
rect 506268 57218 506352 57454
rect 506588 57218 506620 57454
rect 506000 57134 506620 57218
rect 506000 56898 506032 57134
rect 506268 56898 506352 57134
rect 506588 56898 506620 57134
rect 506000 56866 506620 56898
rect 542000 57454 542620 57486
rect 542000 57218 542032 57454
rect 542268 57218 542352 57454
rect 542588 57218 542620 57454
rect 542000 57134 542620 57218
rect 542000 56898 542032 57134
rect 542268 56898 542352 57134
rect 542588 56898 542620 57134
rect 542000 56866 542620 56898
rect 571500 57454 572120 57486
rect 571500 57218 571532 57454
rect 571768 57218 571852 57454
rect 572088 57218 572120 57454
rect 571500 57134 572120 57218
rect 571500 56898 571532 57134
rect 571768 56898 571852 57134
rect 572088 56898 572120 57134
rect 571500 56866 572120 56898
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect 9084 39454 9704 39486
rect 9084 39218 9116 39454
rect 9352 39218 9436 39454
rect 9672 39218 9704 39454
rect 9084 39134 9704 39218
rect 9084 38898 9116 39134
rect 9352 38898 9436 39134
rect 9672 38898 9704 39134
rect 9084 38866 9704 38898
rect 56620 39454 57240 39486
rect 56620 39218 56652 39454
rect 56888 39218 56972 39454
rect 57208 39218 57240 39454
rect 56620 39134 57240 39218
rect 56620 38898 56652 39134
rect 56888 38898 56972 39134
rect 57208 38898 57240 39134
rect 56620 38866 57240 38898
rect 92620 39454 93240 39486
rect 92620 39218 92652 39454
rect 92888 39218 92972 39454
rect 93208 39218 93240 39454
rect 92620 39134 93240 39218
rect 92620 38898 92652 39134
rect 92888 38898 92972 39134
rect 93208 38898 93240 39134
rect 92620 38866 93240 38898
rect 128620 39454 129240 39486
rect 128620 39218 128652 39454
rect 128888 39218 128972 39454
rect 129208 39218 129240 39454
rect 128620 39134 129240 39218
rect 128620 38898 128652 39134
rect 128888 38898 128972 39134
rect 129208 38898 129240 39134
rect 128620 38866 129240 38898
rect 164620 39454 165240 39486
rect 164620 39218 164652 39454
rect 164888 39218 164972 39454
rect 165208 39218 165240 39454
rect 164620 39134 165240 39218
rect 164620 38898 164652 39134
rect 164888 38898 164972 39134
rect 165208 38898 165240 39134
rect 164620 38866 165240 38898
rect 200620 39454 201240 39486
rect 200620 39218 200652 39454
rect 200888 39218 200972 39454
rect 201208 39218 201240 39454
rect 200620 39134 201240 39218
rect 200620 38898 200652 39134
rect 200888 38898 200972 39134
rect 201208 38898 201240 39134
rect 200620 38866 201240 38898
rect 236620 39454 237240 39486
rect 236620 39218 236652 39454
rect 236888 39218 236972 39454
rect 237208 39218 237240 39454
rect 236620 39134 237240 39218
rect 236620 38898 236652 39134
rect 236888 38898 236972 39134
rect 237208 38898 237240 39134
rect 236620 38866 237240 38898
rect 272620 39454 273240 39486
rect 272620 39218 272652 39454
rect 272888 39218 272972 39454
rect 273208 39218 273240 39454
rect 272620 39134 273240 39218
rect 272620 38898 272652 39134
rect 272888 38898 272972 39134
rect 273208 38898 273240 39134
rect 272620 38866 273240 38898
rect 308620 39454 309240 39486
rect 308620 39218 308652 39454
rect 308888 39218 308972 39454
rect 309208 39218 309240 39454
rect 308620 39134 309240 39218
rect 308620 38898 308652 39134
rect 308888 38898 308972 39134
rect 309208 38898 309240 39134
rect 308620 38866 309240 38898
rect 344620 39454 345240 39486
rect 344620 39218 344652 39454
rect 344888 39218 344972 39454
rect 345208 39218 345240 39454
rect 344620 39134 345240 39218
rect 344620 38898 344652 39134
rect 344888 38898 344972 39134
rect 345208 38898 345240 39134
rect 344620 38866 345240 38898
rect 380620 39454 381240 39486
rect 380620 39218 380652 39454
rect 380888 39218 380972 39454
rect 381208 39218 381240 39454
rect 380620 39134 381240 39218
rect 380620 38898 380652 39134
rect 380888 38898 380972 39134
rect 381208 38898 381240 39134
rect 380620 38866 381240 38898
rect 416620 39454 417240 39486
rect 416620 39218 416652 39454
rect 416888 39218 416972 39454
rect 417208 39218 417240 39454
rect 416620 39134 417240 39218
rect 416620 38898 416652 39134
rect 416888 38898 416972 39134
rect 417208 38898 417240 39134
rect 416620 38866 417240 38898
rect 452620 39454 453240 39486
rect 452620 39218 452652 39454
rect 452888 39218 452972 39454
rect 453208 39218 453240 39454
rect 452620 39134 453240 39218
rect 452620 38898 452652 39134
rect 452888 38898 452972 39134
rect 453208 38898 453240 39134
rect 452620 38866 453240 38898
rect 488620 39454 489240 39486
rect 488620 39218 488652 39454
rect 488888 39218 488972 39454
rect 489208 39218 489240 39454
rect 488620 39134 489240 39218
rect 488620 38898 488652 39134
rect 488888 38898 488972 39134
rect 489208 38898 489240 39134
rect 488620 38866 489240 38898
rect 524620 39454 525240 39486
rect 524620 39218 524652 39454
rect 524888 39218 524972 39454
rect 525208 39218 525240 39454
rect 524620 39134 525240 39218
rect 524620 38898 524652 39134
rect 524888 38898 524972 39134
rect 525208 38898 525240 39134
rect 524620 38866 525240 38898
rect 560620 39454 561240 39486
rect 560620 39218 560652 39454
rect 560888 39218 560972 39454
rect 561208 39218 561240 39454
rect 560620 39134 561240 39218
rect 560620 38898 560652 39134
rect 560888 38898 560972 39134
rect 561208 38898 561240 39134
rect 560620 38866 561240 38898
rect 570260 39454 570880 39486
rect 570260 39218 570292 39454
rect 570528 39218 570612 39454
rect 570848 39218 570880 39454
rect 570260 39134 570880 39218
rect 570260 38898 570292 39134
rect 570528 38898 570612 39134
rect 570848 38898 570880 39134
rect 570260 38866 570880 38898
rect 7844 21454 8464 21486
rect 7844 21218 7876 21454
rect 8112 21218 8196 21454
rect 8432 21218 8464 21454
rect 7844 21134 8464 21218
rect 7844 20898 7876 21134
rect 8112 20898 8196 21134
rect 8432 20898 8464 21134
rect 7844 20866 8464 20898
rect 38000 21454 38620 21486
rect 38000 21218 38032 21454
rect 38268 21218 38352 21454
rect 38588 21218 38620 21454
rect 38000 21134 38620 21218
rect 38000 20898 38032 21134
rect 38268 20898 38352 21134
rect 38588 20898 38620 21134
rect 38000 20866 38620 20898
rect 74000 21454 74620 21486
rect 74000 21218 74032 21454
rect 74268 21218 74352 21454
rect 74588 21218 74620 21454
rect 74000 21134 74620 21218
rect 74000 20898 74032 21134
rect 74268 20898 74352 21134
rect 74588 20898 74620 21134
rect 74000 20866 74620 20898
rect 110000 21454 110620 21486
rect 110000 21218 110032 21454
rect 110268 21218 110352 21454
rect 110588 21218 110620 21454
rect 110000 21134 110620 21218
rect 110000 20898 110032 21134
rect 110268 20898 110352 21134
rect 110588 20898 110620 21134
rect 110000 20866 110620 20898
rect 146000 21454 146620 21486
rect 146000 21218 146032 21454
rect 146268 21218 146352 21454
rect 146588 21218 146620 21454
rect 146000 21134 146620 21218
rect 146000 20898 146032 21134
rect 146268 20898 146352 21134
rect 146588 20898 146620 21134
rect 146000 20866 146620 20898
rect 182000 21454 182620 21486
rect 182000 21218 182032 21454
rect 182268 21218 182352 21454
rect 182588 21218 182620 21454
rect 182000 21134 182620 21218
rect 182000 20898 182032 21134
rect 182268 20898 182352 21134
rect 182588 20898 182620 21134
rect 182000 20866 182620 20898
rect 218000 21454 218620 21486
rect 218000 21218 218032 21454
rect 218268 21218 218352 21454
rect 218588 21218 218620 21454
rect 218000 21134 218620 21218
rect 218000 20898 218032 21134
rect 218268 20898 218352 21134
rect 218588 20898 218620 21134
rect 218000 20866 218620 20898
rect 254000 21454 254620 21486
rect 254000 21218 254032 21454
rect 254268 21218 254352 21454
rect 254588 21218 254620 21454
rect 254000 21134 254620 21218
rect 254000 20898 254032 21134
rect 254268 20898 254352 21134
rect 254588 20898 254620 21134
rect 254000 20866 254620 20898
rect 290000 21454 290620 21486
rect 290000 21218 290032 21454
rect 290268 21218 290352 21454
rect 290588 21218 290620 21454
rect 290000 21134 290620 21218
rect 290000 20898 290032 21134
rect 290268 20898 290352 21134
rect 290588 20898 290620 21134
rect 290000 20866 290620 20898
rect 326000 21454 326620 21486
rect 326000 21218 326032 21454
rect 326268 21218 326352 21454
rect 326588 21218 326620 21454
rect 326000 21134 326620 21218
rect 326000 20898 326032 21134
rect 326268 20898 326352 21134
rect 326588 20898 326620 21134
rect 326000 20866 326620 20898
rect 362000 21454 362620 21486
rect 362000 21218 362032 21454
rect 362268 21218 362352 21454
rect 362588 21218 362620 21454
rect 362000 21134 362620 21218
rect 362000 20898 362032 21134
rect 362268 20898 362352 21134
rect 362588 20898 362620 21134
rect 362000 20866 362620 20898
rect 398000 21454 398620 21486
rect 398000 21218 398032 21454
rect 398268 21218 398352 21454
rect 398588 21218 398620 21454
rect 398000 21134 398620 21218
rect 398000 20898 398032 21134
rect 398268 20898 398352 21134
rect 398588 20898 398620 21134
rect 398000 20866 398620 20898
rect 434000 21454 434620 21486
rect 434000 21218 434032 21454
rect 434268 21218 434352 21454
rect 434588 21218 434620 21454
rect 434000 21134 434620 21218
rect 434000 20898 434032 21134
rect 434268 20898 434352 21134
rect 434588 20898 434620 21134
rect 434000 20866 434620 20898
rect 470000 21454 470620 21486
rect 470000 21218 470032 21454
rect 470268 21218 470352 21454
rect 470588 21218 470620 21454
rect 470000 21134 470620 21218
rect 470000 20898 470032 21134
rect 470268 20898 470352 21134
rect 470588 20898 470620 21134
rect 470000 20866 470620 20898
rect 506000 21454 506620 21486
rect 506000 21218 506032 21454
rect 506268 21218 506352 21454
rect 506588 21218 506620 21454
rect 506000 21134 506620 21218
rect 506000 20898 506032 21134
rect 506268 20898 506352 21134
rect 506588 20898 506620 21134
rect 506000 20866 506620 20898
rect 542000 21454 542620 21486
rect 542000 21218 542032 21454
rect 542268 21218 542352 21454
rect 542588 21218 542620 21454
rect 542000 21134 542620 21218
rect 542000 20898 542032 21134
rect 542268 20898 542352 21134
rect 542588 20898 542620 21134
rect 542000 20866 542620 20898
rect 571500 21454 572120 21486
rect 571500 21218 571532 21454
rect 571768 21218 571852 21454
rect 572088 21218 572120 21454
rect 571500 21134 572120 21218
rect 571500 20898 571532 21134
rect 571768 20898 571852 21134
rect 572088 20898 572120 21134
rect 571500 20866 572120 20898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 -346 2414 2000
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 2000
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 2000
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 2000
rect 19794 -1306 20414 2000
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 -3226 24134 2000
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 -5146 27854 2000
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 2000
rect 37794 -346 38414 2000
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 -2266 42134 2000
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 -4186 45854 2000
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 2000
rect 55794 -1306 56414 2000
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 -3226 60134 2000
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 2000
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 2000
rect 73794 -346 74414 2000
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 -2266 78134 2000
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 -4186 81854 2000
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 2000
rect 91794 -1306 92414 2000
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 -3226 96134 2000
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 -5146 99854 2000
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 2000
rect 109794 -346 110414 2000
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 -2266 114134 2000
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 -4186 117854 2000
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 2000
rect 127794 -1306 128414 2000
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 -3226 132134 2000
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 -5146 135854 2000
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 2000
rect 145794 -346 146414 2000
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 -2266 150134 2000
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 -4186 153854 2000
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 2000
rect 163794 -1306 164414 2000
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 -3226 168134 2000
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 2000
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 2000
rect 181794 -346 182414 2000
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 -2266 186134 2000
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 -4186 189854 2000
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 2000
rect 199794 -1306 200414 2000
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 -3226 204134 2000
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 2000
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 2000
rect 217794 -346 218414 2000
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 -2266 222134 2000
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 -4186 225854 2000
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 2000
rect 235794 -1306 236414 2000
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 -3226 240134 2000
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 2000
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 2000
rect 253794 -346 254414 2000
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 -2266 258134 2000
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 -4186 261854 2000
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 2000
rect 271794 -1306 272414 2000
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 -3226 276134 2000
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 2000
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 2000
rect 289794 -346 290414 2000
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 -2266 294134 2000
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 -4186 297854 2000
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 2000
rect 307794 -1306 308414 2000
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 -3226 312134 2000
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 -5146 315854 2000
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 2000
rect 325794 -346 326414 2000
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 -2266 330134 2000
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 -4186 333854 2000
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 2000
rect 343794 -1306 344414 2000
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 -3226 348134 2000
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 -5146 351854 2000
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 2000
rect 361794 -346 362414 2000
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 -2266 366134 2000
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 -4186 369854 2000
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 2000
rect 379794 -1306 380414 2000
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 -3226 384134 2000
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 -5146 387854 2000
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 2000
rect 397794 -346 398414 2000
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 -2266 402134 2000
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 -4186 405854 2000
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 2000
rect 415794 -1306 416414 2000
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 -3226 420134 2000
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 -5146 423854 2000
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 2000
rect 433794 -346 434414 2000
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 -2266 438134 2000
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 -4186 441854 2000
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 2000
rect 451794 -1306 452414 2000
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 -3226 456134 2000
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 -5146 459854 2000
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 2000
rect 469794 -346 470414 2000
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 -2266 474134 2000
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 -4186 477854 2000
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 2000
rect 487794 -1306 488414 2000
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 -3226 492134 2000
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 -5146 495854 2000
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 2000
rect 505794 -346 506414 2000
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 -2266 510134 2000
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 -4186 513854 2000
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 2000
rect 523794 -1306 524414 2000
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 -3226 528134 2000
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 -5146 531854 2000
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 2000
rect 541794 -346 542414 2000
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 -2266 546134 2000
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 -4186 549854 2000
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 2000
rect 559794 -1306 560414 2000
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 -3226 564134 2000
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 -5146 567854 2000
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 2000
rect 577794 -346 578414 2000
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect 9116 687218 9352 687454
rect 9436 687218 9672 687454
rect 9116 686898 9352 687134
rect 9436 686898 9672 687134
rect 56652 687218 56888 687454
rect 56972 687218 57208 687454
rect 56652 686898 56888 687134
rect 56972 686898 57208 687134
rect 92652 687218 92888 687454
rect 92972 687218 93208 687454
rect 92652 686898 92888 687134
rect 92972 686898 93208 687134
rect 128652 687218 128888 687454
rect 128972 687218 129208 687454
rect 128652 686898 128888 687134
rect 128972 686898 129208 687134
rect 164652 687218 164888 687454
rect 164972 687218 165208 687454
rect 164652 686898 164888 687134
rect 164972 686898 165208 687134
rect 200652 687218 200888 687454
rect 200972 687218 201208 687454
rect 200652 686898 200888 687134
rect 200972 686898 201208 687134
rect 236652 687218 236888 687454
rect 236972 687218 237208 687454
rect 236652 686898 236888 687134
rect 236972 686898 237208 687134
rect 272652 687218 272888 687454
rect 272972 687218 273208 687454
rect 272652 686898 272888 687134
rect 272972 686898 273208 687134
rect 308652 687218 308888 687454
rect 308972 687218 309208 687454
rect 308652 686898 308888 687134
rect 308972 686898 309208 687134
rect 344652 687218 344888 687454
rect 344972 687218 345208 687454
rect 344652 686898 344888 687134
rect 344972 686898 345208 687134
rect 380652 687218 380888 687454
rect 380972 687218 381208 687454
rect 380652 686898 380888 687134
rect 380972 686898 381208 687134
rect 416652 687218 416888 687454
rect 416972 687218 417208 687454
rect 416652 686898 416888 687134
rect 416972 686898 417208 687134
rect 452652 687218 452888 687454
rect 452972 687218 453208 687454
rect 452652 686898 452888 687134
rect 452972 686898 453208 687134
rect 488652 687218 488888 687454
rect 488972 687218 489208 687454
rect 488652 686898 488888 687134
rect 488972 686898 489208 687134
rect 524652 687218 524888 687454
rect 524972 687218 525208 687454
rect 524652 686898 524888 687134
rect 524972 686898 525208 687134
rect 560652 687218 560888 687454
rect 560972 687218 561208 687454
rect 560652 686898 560888 687134
rect 560972 686898 561208 687134
rect 570292 687218 570528 687454
rect 570612 687218 570848 687454
rect 570292 686898 570528 687134
rect 570612 686898 570848 687134
rect 7876 669218 8112 669454
rect 8196 669218 8432 669454
rect 7876 668898 8112 669134
rect 8196 668898 8432 669134
rect 38032 669218 38268 669454
rect 38352 669218 38588 669454
rect 38032 668898 38268 669134
rect 38352 668898 38588 669134
rect 74032 669218 74268 669454
rect 74352 669218 74588 669454
rect 74032 668898 74268 669134
rect 74352 668898 74588 669134
rect 100443 669218 100679 669454
rect 100443 668898 100679 669134
rect 198919 669218 199155 669454
rect 198919 668898 199155 669134
rect 216399 669218 216635 669454
rect 216399 668898 216635 669134
rect 314875 669218 315111 669454
rect 314875 668898 315111 669134
rect 326032 669218 326268 669454
rect 326352 669218 326588 669454
rect 326032 668898 326268 669134
rect 326352 668898 326588 669134
rect 332355 669218 332591 669454
rect 332355 668898 332591 669134
rect 430831 669218 431067 669454
rect 430831 668898 431067 669134
rect 434032 669218 434268 669454
rect 434352 669218 434588 669454
rect 434032 668898 434268 669134
rect 434352 668898 434588 669134
rect 448311 669218 448547 669454
rect 448311 668898 448547 669134
rect 546787 669218 547023 669454
rect 546787 668898 547023 669134
rect 571532 669218 571768 669454
rect 571852 669218 572088 669454
rect 571532 668898 571768 669134
rect 571852 668898 572088 669134
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect 9116 651218 9352 651454
rect 9436 651218 9672 651454
rect 9116 650898 9352 651134
rect 9436 650898 9672 651134
rect 56652 651218 56888 651454
rect 56972 651218 57208 651454
rect 56652 650898 56888 651134
rect 56972 650898 57208 651134
rect 92652 651218 92888 651454
rect 92972 651218 93208 651454
rect 92652 650898 92888 651134
rect 92972 650898 93208 651134
rect 101163 651218 101399 651454
rect 101163 650898 101399 651134
rect 198199 651218 198435 651454
rect 198199 650898 198435 651134
rect 200652 651218 200888 651454
rect 200972 651218 201208 651454
rect 200652 650898 200888 651134
rect 200972 650898 201208 651134
rect 217119 651218 217355 651454
rect 217119 650898 217355 651134
rect 314155 651218 314391 651454
rect 314155 650898 314391 651134
rect 333075 651218 333311 651454
rect 333075 650898 333311 651134
rect 430111 651218 430347 651454
rect 430111 650898 430347 651134
rect 449031 651218 449267 651454
rect 449031 650898 449267 651134
rect 546067 651218 546303 651454
rect 546067 650898 546303 651134
rect 560652 651218 560888 651454
rect 560972 651218 561208 651454
rect 560652 650898 560888 651134
rect 560972 650898 561208 651134
rect 570292 651218 570528 651454
rect 570612 651218 570848 651454
rect 570292 650898 570528 651134
rect 570612 650898 570848 651134
rect 7876 633218 8112 633454
rect 8196 633218 8432 633454
rect 7876 632898 8112 633134
rect 8196 632898 8432 633134
rect 38032 633218 38268 633454
rect 38352 633218 38588 633454
rect 38032 632898 38268 633134
rect 38352 632898 38588 633134
rect 74032 633218 74268 633454
rect 74352 633218 74588 633454
rect 74032 632898 74268 633134
rect 74352 632898 74588 633134
rect 100443 633218 100679 633454
rect 100443 632898 100679 633134
rect 198919 633218 199155 633454
rect 198919 632898 199155 633134
rect 216399 633218 216635 633454
rect 216399 632898 216635 633134
rect 314875 633218 315111 633454
rect 314875 632898 315111 633134
rect 326032 633218 326268 633454
rect 326352 633218 326588 633454
rect 326032 632898 326268 633134
rect 326352 632898 326588 633134
rect 332355 633218 332591 633454
rect 332355 632898 332591 633134
rect 430831 633218 431067 633454
rect 430831 632898 431067 633134
rect 434032 633218 434268 633454
rect 434352 633218 434588 633454
rect 434032 632898 434268 633134
rect 434352 632898 434588 633134
rect 448311 633218 448547 633454
rect 448311 632898 448547 633134
rect 546787 633218 547023 633454
rect 546787 632898 547023 633134
rect 571532 633218 571768 633454
rect 571852 633218 572088 633454
rect 571532 632898 571768 633134
rect 571852 632898 572088 633134
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect 9116 615218 9352 615454
rect 9436 615218 9672 615454
rect 9116 614898 9352 615134
rect 9436 614898 9672 615134
rect 56652 615218 56888 615454
rect 56972 615218 57208 615454
rect 56652 614898 56888 615134
rect 56972 614898 57208 615134
rect 92652 615218 92888 615454
rect 92972 615218 93208 615454
rect 92652 614898 92888 615134
rect 92972 614898 93208 615134
rect 101163 615218 101399 615454
rect 101163 614898 101399 615134
rect 198199 615218 198435 615454
rect 198199 614898 198435 615134
rect 200652 615218 200888 615454
rect 200972 615218 201208 615454
rect 200652 614898 200888 615134
rect 200972 614898 201208 615134
rect 217119 615218 217355 615454
rect 217119 614898 217355 615134
rect 314155 615218 314391 615454
rect 314155 614898 314391 615134
rect 333075 615218 333311 615454
rect 333075 614898 333311 615134
rect 430111 615218 430347 615454
rect 430111 614898 430347 615134
rect 449031 615218 449267 615454
rect 449031 614898 449267 615134
rect 546067 615218 546303 615454
rect 546067 614898 546303 615134
rect 560652 615218 560888 615454
rect 560972 615218 561208 615454
rect 560652 614898 560888 615134
rect 560972 614898 561208 615134
rect 570292 615218 570528 615454
rect 570612 615218 570848 615454
rect 570292 614898 570528 615134
rect 570612 614898 570848 615134
rect 7876 597218 8112 597454
rect 8196 597218 8432 597454
rect 7876 596898 8112 597134
rect 8196 596898 8432 597134
rect 38032 597218 38268 597454
rect 38352 597218 38588 597454
rect 38032 596898 38268 597134
rect 38352 596898 38588 597134
rect 74032 597218 74268 597454
rect 74352 597218 74588 597454
rect 74032 596898 74268 597134
rect 74352 596898 74588 597134
rect 100443 597218 100679 597454
rect 100443 596898 100679 597134
rect 198919 597218 199155 597454
rect 198919 596898 199155 597134
rect 216399 597218 216635 597454
rect 216399 596898 216635 597134
rect 314875 597218 315111 597454
rect 314875 596898 315111 597134
rect 326032 597218 326268 597454
rect 326352 597218 326588 597454
rect 326032 596898 326268 597134
rect 326352 596898 326588 597134
rect 332355 597218 332591 597454
rect 332355 596898 332591 597134
rect 430831 597218 431067 597454
rect 430831 596898 431067 597134
rect 434032 597218 434268 597454
rect 434352 597218 434588 597454
rect 434032 596898 434268 597134
rect 434352 596898 434588 597134
rect 448311 597218 448547 597454
rect 448311 596898 448547 597134
rect 546787 597218 547023 597454
rect 546787 596898 547023 597134
rect 571532 597218 571768 597454
rect 571852 597218 572088 597454
rect 571532 596898 571768 597134
rect 571852 596898 572088 597134
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect 9116 579218 9352 579454
rect 9436 579218 9672 579454
rect 9116 578898 9352 579134
rect 9436 578898 9672 579134
rect 56652 579218 56888 579454
rect 56972 579218 57208 579454
rect 56652 578898 56888 579134
rect 56972 578898 57208 579134
rect 92652 579218 92888 579454
rect 92972 579218 93208 579454
rect 92652 578898 92888 579134
rect 92972 578898 93208 579134
rect 128652 579218 128888 579454
rect 128972 579218 129208 579454
rect 128652 578898 128888 579134
rect 128972 578898 129208 579134
rect 164652 579218 164888 579454
rect 164972 579218 165208 579454
rect 164652 578898 164888 579134
rect 164972 578898 165208 579134
rect 200652 579218 200888 579454
rect 200972 579218 201208 579454
rect 200652 578898 200888 579134
rect 200972 578898 201208 579134
rect 236652 579218 236888 579454
rect 236972 579218 237208 579454
rect 236652 578898 236888 579134
rect 236972 578898 237208 579134
rect 272652 579218 272888 579454
rect 272972 579218 273208 579454
rect 272652 578898 272888 579134
rect 272972 578898 273208 579134
rect 308652 579218 308888 579454
rect 308972 579218 309208 579454
rect 308652 578898 308888 579134
rect 308972 578898 309208 579134
rect 344652 579218 344888 579454
rect 344972 579218 345208 579454
rect 344652 578898 344888 579134
rect 344972 578898 345208 579134
rect 380652 579218 380888 579454
rect 380972 579218 381208 579454
rect 380652 578898 380888 579134
rect 380972 578898 381208 579134
rect 416652 579218 416888 579454
rect 416972 579218 417208 579454
rect 416652 578898 416888 579134
rect 416972 578898 417208 579134
rect 452652 579218 452888 579454
rect 452972 579218 453208 579454
rect 452652 578898 452888 579134
rect 452972 578898 453208 579134
rect 488652 579218 488888 579454
rect 488972 579218 489208 579454
rect 488652 578898 488888 579134
rect 488972 578898 489208 579134
rect 524652 579218 524888 579454
rect 524972 579218 525208 579454
rect 524652 578898 524888 579134
rect 524972 578898 525208 579134
rect 560652 579218 560888 579454
rect 560972 579218 561208 579454
rect 560652 578898 560888 579134
rect 560972 578898 561208 579134
rect 570292 579218 570528 579454
rect 570612 579218 570848 579454
rect 570292 578898 570528 579134
rect 570612 578898 570848 579134
rect 7876 561218 8112 561454
rect 8196 561218 8432 561454
rect 7876 560898 8112 561134
rect 8196 560898 8432 561134
rect 38032 561218 38268 561454
rect 38352 561218 38588 561454
rect 38032 560898 38268 561134
rect 38352 560898 38588 561134
rect 74032 561218 74268 561454
rect 74352 561218 74588 561454
rect 74032 560898 74268 561134
rect 74352 560898 74588 561134
rect 110032 561218 110268 561454
rect 110352 561218 110588 561454
rect 110032 560898 110268 561134
rect 110352 560898 110588 561134
rect 146032 561218 146268 561454
rect 146352 561218 146588 561454
rect 146032 560898 146268 561134
rect 146352 560898 146588 561134
rect 182032 561218 182268 561454
rect 182352 561218 182588 561454
rect 182032 560898 182268 561134
rect 182352 560898 182588 561134
rect 218032 561218 218268 561454
rect 218352 561218 218588 561454
rect 218032 560898 218268 561134
rect 218352 560898 218588 561134
rect 254032 561218 254268 561454
rect 254352 561218 254588 561454
rect 254032 560898 254268 561134
rect 254352 560898 254588 561134
rect 290032 561218 290268 561454
rect 290352 561218 290588 561454
rect 290032 560898 290268 561134
rect 290352 560898 290588 561134
rect 326032 561218 326268 561454
rect 326352 561218 326588 561454
rect 326032 560898 326268 561134
rect 326352 560898 326588 561134
rect 332355 561218 332591 561454
rect 332355 560898 332591 561134
rect 430831 561218 431067 561454
rect 430831 560898 431067 561134
rect 434032 561218 434268 561454
rect 434352 561218 434588 561454
rect 434032 560898 434268 561134
rect 434352 560898 434588 561134
rect 448311 561218 448547 561454
rect 448311 560898 448547 561134
rect 546787 561218 547023 561454
rect 546787 560898 547023 561134
rect 571532 561218 571768 561454
rect 571852 561218 572088 561454
rect 571532 560898 571768 561134
rect 571852 560898 572088 561134
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect 9116 543218 9352 543454
rect 9436 543218 9672 543454
rect 9116 542898 9352 543134
rect 9436 542898 9672 543134
rect 56652 543218 56888 543454
rect 56972 543218 57208 543454
rect 56652 542898 56888 543134
rect 56972 542898 57208 543134
rect 92652 543218 92888 543454
rect 92972 543218 93208 543454
rect 92652 542898 92888 543134
rect 92972 542898 93208 543134
rect 128652 543218 128888 543454
rect 128972 543218 129208 543454
rect 128652 542898 128888 543134
rect 128972 542898 129208 543134
rect 164652 543218 164888 543454
rect 164972 543218 165208 543454
rect 164652 542898 164888 543134
rect 164972 542898 165208 543134
rect 200652 543218 200888 543454
rect 200972 543218 201208 543454
rect 200652 542898 200888 543134
rect 200972 542898 201208 543134
rect 236652 543218 236888 543454
rect 236972 543218 237208 543454
rect 236652 542898 236888 543134
rect 236972 542898 237208 543134
rect 272652 543218 272888 543454
rect 272972 543218 273208 543454
rect 272652 542898 272888 543134
rect 272972 542898 273208 543134
rect 308652 543218 308888 543454
rect 308972 543218 309208 543454
rect 308652 542898 308888 543134
rect 308972 542898 309208 543134
rect 333075 543218 333311 543454
rect 333075 542898 333311 543134
rect 430111 543218 430347 543454
rect 430111 542898 430347 543134
rect 449031 543218 449267 543454
rect 449031 542898 449267 543134
rect 546067 543218 546303 543454
rect 546067 542898 546303 543134
rect 560652 543218 560888 543454
rect 560972 543218 561208 543454
rect 560652 542898 560888 543134
rect 560972 542898 561208 543134
rect 570292 543218 570528 543454
rect 570612 543218 570848 543454
rect 570292 542898 570528 543134
rect 570612 542898 570848 543134
rect 7876 525218 8112 525454
rect 8196 525218 8432 525454
rect 7876 524898 8112 525134
rect 8196 524898 8432 525134
rect 38032 525218 38268 525454
rect 38352 525218 38588 525454
rect 38032 524898 38268 525134
rect 38352 524898 38588 525134
rect 74032 525218 74268 525454
rect 74352 525218 74588 525454
rect 74032 524898 74268 525134
rect 74352 524898 74588 525134
rect 110032 525218 110268 525454
rect 110352 525218 110588 525454
rect 110032 524898 110268 525134
rect 110352 524898 110588 525134
rect 146032 525218 146268 525454
rect 146352 525218 146588 525454
rect 146032 524898 146268 525134
rect 146352 524898 146588 525134
rect 182032 525218 182268 525454
rect 182352 525218 182588 525454
rect 182032 524898 182268 525134
rect 182352 524898 182588 525134
rect 218032 525218 218268 525454
rect 218352 525218 218588 525454
rect 218032 524898 218268 525134
rect 218352 524898 218588 525134
rect 254032 525218 254268 525454
rect 254352 525218 254588 525454
rect 254032 524898 254268 525134
rect 254352 524898 254588 525134
rect 290032 525218 290268 525454
rect 290352 525218 290588 525454
rect 290032 524898 290268 525134
rect 290352 524898 290588 525134
rect 326032 525218 326268 525454
rect 326352 525218 326588 525454
rect 326032 524898 326268 525134
rect 326352 524898 326588 525134
rect 332355 525218 332591 525454
rect 332355 524898 332591 525134
rect 430831 525218 431067 525454
rect 430831 524898 431067 525134
rect 434032 525218 434268 525454
rect 434352 525218 434588 525454
rect 434032 524898 434268 525134
rect 434352 524898 434588 525134
rect 448311 525218 448547 525454
rect 448311 524898 448547 525134
rect 546787 525218 547023 525454
rect 546787 524898 547023 525134
rect 571532 525218 571768 525454
rect 571852 525218 572088 525454
rect 571532 524898 571768 525134
rect 571852 524898 572088 525134
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect 9116 507218 9352 507454
rect 9436 507218 9672 507454
rect 9116 506898 9352 507134
rect 9436 506898 9672 507134
rect 56652 507218 56888 507454
rect 56972 507218 57208 507454
rect 56652 506898 56888 507134
rect 56972 506898 57208 507134
rect 92652 507218 92888 507454
rect 92972 507218 93208 507454
rect 92652 506898 92888 507134
rect 92972 506898 93208 507134
rect 128652 507218 128888 507454
rect 128972 507218 129208 507454
rect 128652 506898 128888 507134
rect 128972 506898 129208 507134
rect 164652 507218 164888 507454
rect 164972 507218 165208 507454
rect 164652 506898 164888 507134
rect 164972 506898 165208 507134
rect 200652 507218 200888 507454
rect 200972 507218 201208 507454
rect 200652 506898 200888 507134
rect 200972 506898 201208 507134
rect 236652 507218 236888 507454
rect 236972 507218 237208 507454
rect 236652 506898 236888 507134
rect 236972 506898 237208 507134
rect 272652 507218 272888 507454
rect 272972 507218 273208 507454
rect 272652 506898 272888 507134
rect 272972 506898 273208 507134
rect 308652 507218 308888 507454
rect 308972 507218 309208 507454
rect 308652 506898 308888 507134
rect 308972 506898 309208 507134
rect 333075 507218 333311 507454
rect 333075 506898 333311 507134
rect 430111 507218 430347 507454
rect 430111 506898 430347 507134
rect 449031 507218 449267 507454
rect 449031 506898 449267 507134
rect 546067 507218 546303 507454
rect 546067 506898 546303 507134
rect 560652 507218 560888 507454
rect 560972 507218 561208 507454
rect 560652 506898 560888 507134
rect 560972 506898 561208 507134
rect 570292 507218 570528 507454
rect 570612 507218 570848 507454
rect 570292 506898 570528 507134
rect 570612 506898 570848 507134
rect 7876 489218 8112 489454
rect 8196 489218 8432 489454
rect 7876 488898 8112 489134
rect 8196 488898 8432 489134
rect 38032 489218 38268 489454
rect 38352 489218 38588 489454
rect 38032 488898 38268 489134
rect 38352 488898 38588 489134
rect 74032 489218 74268 489454
rect 74352 489218 74588 489454
rect 74032 488898 74268 489134
rect 74352 488898 74588 489134
rect 110032 489218 110268 489454
rect 110352 489218 110588 489454
rect 110032 488898 110268 489134
rect 110352 488898 110588 489134
rect 146032 489218 146268 489454
rect 146352 489218 146588 489454
rect 146032 488898 146268 489134
rect 146352 488898 146588 489134
rect 182032 489218 182268 489454
rect 182352 489218 182588 489454
rect 182032 488898 182268 489134
rect 182352 488898 182588 489134
rect 218032 489218 218268 489454
rect 218352 489218 218588 489454
rect 218032 488898 218268 489134
rect 218352 488898 218588 489134
rect 254032 489218 254268 489454
rect 254352 489218 254588 489454
rect 254032 488898 254268 489134
rect 254352 488898 254588 489134
rect 290032 489218 290268 489454
rect 290352 489218 290588 489454
rect 290032 488898 290268 489134
rect 290352 488898 290588 489134
rect 326032 489218 326268 489454
rect 326352 489218 326588 489454
rect 326032 488898 326268 489134
rect 326352 488898 326588 489134
rect 362032 489218 362268 489454
rect 362352 489218 362588 489454
rect 362032 488898 362268 489134
rect 362352 488898 362588 489134
rect 398032 489218 398268 489454
rect 398352 489218 398588 489454
rect 398032 488898 398268 489134
rect 398352 488898 398588 489134
rect 434032 489218 434268 489454
rect 434352 489218 434588 489454
rect 434032 488898 434268 489134
rect 434352 488898 434588 489134
rect 470032 489218 470268 489454
rect 470352 489218 470588 489454
rect 470032 488898 470268 489134
rect 470352 488898 470588 489134
rect 506032 489218 506268 489454
rect 506352 489218 506588 489454
rect 506032 488898 506268 489134
rect 506352 488898 506588 489134
rect 542032 489218 542268 489454
rect 542352 489218 542588 489454
rect 542032 488898 542268 489134
rect 542352 488898 542588 489134
rect 571532 489218 571768 489454
rect 571852 489218 572088 489454
rect 571532 488898 571768 489134
rect 571852 488898 572088 489134
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect 9116 471218 9352 471454
rect 9436 471218 9672 471454
rect 9116 470898 9352 471134
rect 9436 470898 9672 471134
rect 56652 471218 56888 471454
rect 56972 471218 57208 471454
rect 56652 470898 56888 471134
rect 56972 470898 57208 471134
rect 92652 471218 92888 471454
rect 92972 471218 93208 471454
rect 92652 470898 92888 471134
rect 92972 470898 93208 471134
rect 128652 471218 128888 471454
rect 128972 471218 129208 471454
rect 128652 470898 128888 471134
rect 128972 470898 129208 471134
rect 164652 471218 164888 471454
rect 164972 471218 165208 471454
rect 164652 470898 164888 471134
rect 164972 470898 165208 471134
rect 200652 471218 200888 471454
rect 200972 471218 201208 471454
rect 200652 470898 200888 471134
rect 200972 470898 201208 471134
rect 236652 471218 236888 471454
rect 236972 471218 237208 471454
rect 236652 470898 236888 471134
rect 236972 470898 237208 471134
rect 272652 471218 272888 471454
rect 272972 471218 273208 471454
rect 272652 470898 272888 471134
rect 272972 470898 273208 471134
rect 308652 471218 308888 471454
rect 308972 471218 309208 471454
rect 308652 470898 308888 471134
rect 308972 470898 309208 471134
rect 333075 471218 333311 471454
rect 333075 470898 333311 471134
rect 430111 471218 430347 471454
rect 430111 470898 430347 471134
rect 449031 471218 449267 471454
rect 449031 470898 449267 471134
rect 546067 471218 546303 471454
rect 546067 470898 546303 471134
rect 560652 471218 560888 471454
rect 560972 471218 561208 471454
rect 560652 470898 560888 471134
rect 560972 470898 561208 471134
rect 570292 471218 570528 471454
rect 570612 471218 570848 471454
rect 570292 470898 570528 471134
rect 570612 470898 570848 471134
rect 7876 453218 8112 453454
rect 8196 453218 8432 453454
rect 7876 452898 8112 453134
rect 8196 452898 8432 453134
rect 38032 453218 38268 453454
rect 38352 453218 38588 453454
rect 38032 452898 38268 453134
rect 38352 452898 38588 453134
rect 74032 453218 74268 453454
rect 74352 453218 74588 453454
rect 74032 452898 74268 453134
rect 74352 452898 74588 453134
rect 110032 453218 110268 453454
rect 110352 453218 110588 453454
rect 110032 452898 110268 453134
rect 110352 452898 110588 453134
rect 146032 453218 146268 453454
rect 146352 453218 146588 453454
rect 146032 452898 146268 453134
rect 146352 452898 146588 453134
rect 182032 453218 182268 453454
rect 182352 453218 182588 453454
rect 182032 452898 182268 453134
rect 182352 452898 182588 453134
rect 218032 453218 218268 453454
rect 218352 453218 218588 453454
rect 218032 452898 218268 453134
rect 218352 452898 218588 453134
rect 254032 453218 254268 453454
rect 254352 453218 254588 453454
rect 254032 452898 254268 453134
rect 254352 452898 254588 453134
rect 290032 453218 290268 453454
rect 290352 453218 290588 453454
rect 290032 452898 290268 453134
rect 290352 452898 290588 453134
rect 326032 453218 326268 453454
rect 326352 453218 326588 453454
rect 326032 452898 326268 453134
rect 326352 452898 326588 453134
rect 332355 453218 332591 453454
rect 332355 452898 332591 453134
rect 430831 453218 431067 453454
rect 430831 452898 431067 453134
rect 434032 453218 434268 453454
rect 434352 453218 434588 453454
rect 434032 452898 434268 453134
rect 434352 452898 434588 453134
rect 448311 453218 448547 453454
rect 448311 452898 448547 453134
rect 546787 453218 547023 453454
rect 546787 452898 547023 453134
rect 571532 453218 571768 453454
rect 571852 453218 572088 453454
rect 571532 452898 571768 453134
rect 571852 452898 572088 453134
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect 9116 435218 9352 435454
rect 9436 435218 9672 435454
rect 9116 434898 9352 435134
rect 9436 434898 9672 435134
rect 56652 435218 56888 435454
rect 56972 435218 57208 435454
rect 56652 434898 56888 435134
rect 56972 434898 57208 435134
rect 92652 435218 92888 435454
rect 92972 435218 93208 435454
rect 92652 434898 92888 435134
rect 92972 434898 93208 435134
rect 128652 435218 128888 435454
rect 128972 435218 129208 435454
rect 128652 434898 128888 435134
rect 128972 434898 129208 435134
rect 164652 435218 164888 435454
rect 164972 435218 165208 435454
rect 164652 434898 164888 435134
rect 164972 434898 165208 435134
rect 200652 435218 200888 435454
rect 200972 435218 201208 435454
rect 200652 434898 200888 435134
rect 200972 434898 201208 435134
rect 236652 435218 236888 435454
rect 236972 435218 237208 435454
rect 236652 434898 236888 435134
rect 236972 434898 237208 435134
rect 272652 435218 272888 435454
rect 272972 435218 273208 435454
rect 272652 434898 272888 435134
rect 272972 434898 273208 435134
rect 308652 435218 308888 435454
rect 308972 435218 309208 435454
rect 308652 434898 308888 435134
rect 308972 434898 309208 435134
rect 333075 435218 333311 435454
rect 333075 434898 333311 435134
rect 430111 435218 430347 435454
rect 430111 434898 430347 435134
rect 449031 435218 449267 435454
rect 449031 434898 449267 435134
rect 546067 435218 546303 435454
rect 546067 434898 546303 435134
rect 560652 435218 560888 435454
rect 560972 435218 561208 435454
rect 560652 434898 560888 435134
rect 560972 434898 561208 435134
rect 570292 435218 570528 435454
rect 570612 435218 570848 435454
rect 570292 434898 570528 435134
rect 570612 434898 570848 435134
rect 7876 417218 8112 417454
rect 8196 417218 8432 417454
rect 7876 416898 8112 417134
rect 8196 416898 8432 417134
rect 38032 417218 38268 417454
rect 38352 417218 38588 417454
rect 38032 416898 38268 417134
rect 38352 416898 38588 417134
rect 74032 417218 74268 417454
rect 74352 417218 74588 417454
rect 74032 416898 74268 417134
rect 74352 416898 74588 417134
rect 110032 417218 110268 417454
rect 110352 417218 110588 417454
rect 110032 416898 110268 417134
rect 110352 416898 110588 417134
rect 146032 417218 146268 417454
rect 146352 417218 146588 417454
rect 146032 416898 146268 417134
rect 146352 416898 146588 417134
rect 182032 417218 182268 417454
rect 182352 417218 182588 417454
rect 182032 416898 182268 417134
rect 182352 416898 182588 417134
rect 218032 417218 218268 417454
rect 218352 417218 218588 417454
rect 218032 416898 218268 417134
rect 218352 416898 218588 417134
rect 254032 417218 254268 417454
rect 254352 417218 254588 417454
rect 254032 416898 254268 417134
rect 254352 416898 254588 417134
rect 290032 417218 290268 417454
rect 290352 417218 290588 417454
rect 290032 416898 290268 417134
rect 290352 416898 290588 417134
rect 326032 417218 326268 417454
rect 326352 417218 326588 417454
rect 326032 416898 326268 417134
rect 326352 416898 326588 417134
rect 332355 417218 332591 417454
rect 332355 416898 332591 417134
rect 430831 417218 431067 417454
rect 430831 416898 431067 417134
rect 434032 417218 434268 417454
rect 434352 417218 434588 417454
rect 434032 416898 434268 417134
rect 434352 416898 434588 417134
rect 448311 417218 448547 417454
rect 448311 416898 448547 417134
rect 546787 417218 547023 417454
rect 546787 416898 547023 417134
rect 571532 417218 571768 417454
rect 571852 417218 572088 417454
rect 571532 416898 571768 417134
rect 571852 416898 572088 417134
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect 9116 399218 9352 399454
rect 9436 399218 9672 399454
rect 9116 398898 9352 399134
rect 9436 398898 9672 399134
rect 56652 399218 56888 399454
rect 56972 399218 57208 399454
rect 56652 398898 56888 399134
rect 56972 398898 57208 399134
rect 92652 399218 92888 399454
rect 92972 399218 93208 399454
rect 92652 398898 92888 399134
rect 92972 398898 93208 399134
rect 128652 399218 128888 399454
rect 128972 399218 129208 399454
rect 128652 398898 128888 399134
rect 128972 398898 129208 399134
rect 164652 399218 164888 399454
rect 164972 399218 165208 399454
rect 164652 398898 164888 399134
rect 164972 398898 165208 399134
rect 200652 399218 200888 399454
rect 200972 399218 201208 399454
rect 200652 398898 200888 399134
rect 200972 398898 201208 399134
rect 236652 399218 236888 399454
rect 236972 399218 237208 399454
rect 236652 398898 236888 399134
rect 236972 398898 237208 399134
rect 272652 399218 272888 399454
rect 272972 399218 273208 399454
rect 272652 398898 272888 399134
rect 272972 398898 273208 399134
rect 308652 399218 308888 399454
rect 308972 399218 309208 399454
rect 308652 398898 308888 399134
rect 308972 398898 309208 399134
rect 333075 399218 333311 399454
rect 333075 398898 333311 399134
rect 430111 399218 430347 399454
rect 430111 398898 430347 399134
rect 449031 399218 449267 399454
rect 449031 398898 449267 399134
rect 546067 399218 546303 399454
rect 546067 398898 546303 399134
rect 560652 399218 560888 399454
rect 560972 399218 561208 399454
rect 560652 398898 560888 399134
rect 560972 398898 561208 399134
rect 570292 399218 570528 399454
rect 570612 399218 570848 399454
rect 570292 398898 570528 399134
rect 570612 398898 570848 399134
rect 7876 381218 8112 381454
rect 8196 381218 8432 381454
rect 7876 380898 8112 381134
rect 8196 380898 8432 381134
rect 38032 381218 38268 381454
rect 38352 381218 38588 381454
rect 38032 380898 38268 381134
rect 38352 380898 38588 381134
rect 74032 381218 74268 381454
rect 74352 381218 74588 381454
rect 74032 380898 74268 381134
rect 74352 380898 74588 381134
rect 110032 381218 110268 381454
rect 110352 381218 110588 381454
rect 110032 380898 110268 381134
rect 110352 380898 110588 381134
rect 146032 381218 146268 381454
rect 146352 381218 146588 381454
rect 146032 380898 146268 381134
rect 146352 380898 146588 381134
rect 182032 381218 182268 381454
rect 182352 381218 182588 381454
rect 182032 380898 182268 381134
rect 182352 380898 182588 381134
rect 218032 381218 218268 381454
rect 218352 381218 218588 381454
rect 218032 380898 218268 381134
rect 218352 380898 218588 381134
rect 254032 381218 254268 381454
rect 254352 381218 254588 381454
rect 254032 380898 254268 381134
rect 254352 380898 254588 381134
rect 290032 381218 290268 381454
rect 290352 381218 290588 381454
rect 290032 380898 290268 381134
rect 290352 380898 290588 381134
rect 326032 381218 326268 381454
rect 326352 381218 326588 381454
rect 326032 380898 326268 381134
rect 326352 380898 326588 381134
rect 362032 381218 362268 381454
rect 362352 381218 362588 381454
rect 362032 380898 362268 381134
rect 362352 380898 362588 381134
rect 398032 381218 398268 381454
rect 398352 381218 398588 381454
rect 398032 380898 398268 381134
rect 398352 380898 398588 381134
rect 434032 381218 434268 381454
rect 434352 381218 434588 381454
rect 434032 380898 434268 381134
rect 434352 380898 434588 381134
rect 470032 381218 470268 381454
rect 470352 381218 470588 381454
rect 470032 380898 470268 381134
rect 470352 380898 470588 381134
rect 506032 381218 506268 381454
rect 506352 381218 506588 381454
rect 506032 380898 506268 381134
rect 506352 380898 506588 381134
rect 542032 381218 542268 381454
rect 542352 381218 542588 381454
rect 542032 380898 542268 381134
rect 542352 380898 542588 381134
rect 571532 381218 571768 381454
rect 571852 381218 572088 381454
rect 571532 380898 571768 381134
rect 571852 380898 572088 381134
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect 9116 363218 9352 363454
rect 9436 363218 9672 363454
rect 9116 362898 9352 363134
rect 9436 362898 9672 363134
rect 56652 363218 56888 363454
rect 56972 363218 57208 363454
rect 56652 362898 56888 363134
rect 56972 362898 57208 363134
rect 92652 363218 92888 363454
rect 92972 363218 93208 363454
rect 92652 362898 92888 363134
rect 92972 362898 93208 363134
rect 128652 363218 128888 363454
rect 128972 363218 129208 363454
rect 128652 362898 128888 363134
rect 128972 362898 129208 363134
rect 164652 363218 164888 363454
rect 164972 363218 165208 363454
rect 164652 362898 164888 363134
rect 164972 362898 165208 363134
rect 200652 363218 200888 363454
rect 200972 363218 201208 363454
rect 200652 362898 200888 363134
rect 200972 362898 201208 363134
rect 236652 363218 236888 363454
rect 236972 363218 237208 363454
rect 236652 362898 236888 363134
rect 236972 362898 237208 363134
rect 272652 363218 272888 363454
rect 272972 363218 273208 363454
rect 272652 362898 272888 363134
rect 272972 362898 273208 363134
rect 308652 363218 308888 363454
rect 308972 363218 309208 363454
rect 308652 362898 308888 363134
rect 308972 362898 309208 363134
rect 333075 363218 333311 363454
rect 333075 362898 333311 363134
rect 430111 363218 430347 363454
rect 430111 362898 430347 363134
rect 449031 363218 449267 363454
rect 449031 362898 449267 363134
rect 546067 363218 546303 363454
rect 546067 362898 546303 363134
rect 560652 363218 560888 363454
rect 560972 363218 561208 363454
rect 560652 362898 560888 363134
rect 560972 362898 561208 363134
rect 570292 363218 570528 363454
rect 570612 363218 570848 363454
rect 570292 362898 570528 363134
rect 570612 362898 570848 363134
rect 7876 345218 8112 345454
rect 8196 345218 8432 345454
rect 7876 344898 8112 345134
rect 8196 344898 8432 345134
rect 38032 345218 38268 345454
rect 38352 345218 38588 345454
rect 38032 344898 38268 345134
rect 38352 344898 38588 345134
rect 74032 345218 74268 345454
rect 74352 345218 74588 345454
rect 74032 344898 74268 345134
rect 74352 344898 74588 345134
rect 110032 345218 110268 345454
rect 110352 345218 110588 345454
rect 110032 344898 110268 345134
rect 110352 344898 110588 345134
rect 146032 345218 146268 345454
rect 146352 345218 146588 345454
rect 146032 344898 146268 345134
rect 146352 344898 146588 345134
rect 182032 345218 182268 345454
rect 182352 345218 182588 345454
rect 182032 344898 182268 345134
rect 182352 344898 182588 345134
rect 218032 345218 218268 345454
rect 218352 345218 218588 345454
rect 218032 344898 218268 345134
rect 218352 344898 218588 345134
rect 254032 345218 254268 345454
rect 254352 345218 254588 345454
rect 254032 344898 254268 345134
rect 254352 344898 254588 345134
rect 290032 345218 290268 345454
rect 290352 345218 290588 345454
rect 290032 344898 290268 345134
rect 290352 344898 290588 345134
rect 326032 345218 326268 345454
rect 326352 345218 326588 345454
rect 326032 344898 326268 345134
rect 326352 344898 326588 345134
rect 332355 345218 332591 345454
rect 332355 344898 332591 345134
rect 430831 345218 431067 345454
rect 430831 344898 431067 345134
rect 434032 345218 434268 345454
rect 434352 345218 434588 345454
rect 434032 344898 434268 345134
rect 434352 344898 434588 345134
rect 448311 345218 448547 345454
rect 448311 344898 448547 345134
rect 546787 345218 547023 345454
rect 546787 344898 547023 345134
rect 571532 345218 571768 345454
rect 571852 345218 572088 345454
rect 571532 344898 571768 345134
rect 571852 344898 572088 345134
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect 9116 327218 9352 327454
rect 9436 327218 9672 327454
rect 9116 326898 9352 327134
rect 9436 326898 9672 327134
rect 56652 327218 56888 327454
rect 56972 327218 57208 327454
rect 56652 326898 56888 327134
rect 56972 326898 57208 327134
rect 92652 327218 92888 327454
rect 92972 327218 93208 327454
rect 92652 326898 92888 327134
rect 92972 326898 93208 327134
rect 128652 327218 128888 327454
rect 128972 327218 129208 327454
rect 128652 326898 128888 327134
rect 128972 326898 129208 327134
rect 164652 327218 164888 327454
rect 164972 327218 165208 327454
rect 164652 326898 164888 327134
rect 164972 326898 165208 327134
rect 200652 327218 200888 327454
rect 200972 327218 201208 327454
rect 200652 326898 200888 327134
rect 200972 326898 201208 327134
rect 236652 327218 236888 327454
rect 236972 327218 237208 327454
rect 236652 326898 236888 327134
rect 236972 326898 237208 327134
rect 272652 327218 272888 327454
rect 272972 327218 273208 327454
rect 272652 326898 272888 327134
rect 272972 326898 273208 327134
rect 308652 327218 308888 327454
rect 308972 327218 309208 327454
rect 308652 326898 308888 327134
rect 308972 326898 309208 327134
rect 333075 327218 333311 327454
rect 333075 326898 333311 327134
rect 430111 327218 430347 327454
rect 430111 326898 430347 327134
rect 449031 327218 449267 327454
rect 449031 326898 449267 327134
rect 546067 327218 546303 327454
rect 546067 326898 546303 327134
rect 560652 327218 560888 327454
rect 560972 327218 561208 327454
rect 560652 326898 560888 327134
rect 560972 326898 561208 327134
rect 570292 327218 570528 327454
rect 570612 327218 570848 327454
rect 570292 326898 570528 327134
rect 570612 326898 570848 327134
rect 7876 309218 8112 309454
rect 8196 309218 8432 309454
rect 7876 308898 8112 309134
rect 8196 308898 8432 309134
rect 38032 309218 38268 309454
rect 38352 309218 38588 309454
rect 38032 308898 38268 309134
rect 38352 308898 38588 309134
rect 74032 309218 74268 309454
rect 74352 309218 74588 309454
rect 74032 308898 74268 309134
rect 74352 308898 74588 309134
rect 110032 309218 110268 309454
rect 110352 309218 110588 309454
rect 110032 308898 110268 309134
rect 110352 308898 110588 309134
rect 146032 309218 146268 309454
rect 146352 309218 146588 309454
rect 146032 308898 146268 309134
rect 146352 308898 146588 309134
rect 182032 309218 182268 309454
rect 182352 309218 182588 309454
rect 182032 308898 182268 309134
rect 182352 308898 182588 309134
rect 218032 309218 218268 309454
rect 218352 309218 218588 309454
rect 218032 308898 218268 309134
rect 218352 308898 218588 309134
rect 254032 309218 254268 309454
rect 254352 309218 254588 309454
rect 254032 308898 254268 309134
rect 254352 308898 254588 309134
rect 290032 309218 290268 309454
rect 290352 309218 290588 309454
rect 290032 308898 290268 309134
rect 290352 308898 290588 309134
rect 326032 309218 326268 309454
rect 326352 309218 326588 309454
rect 326032 308898 326268 309134
rect 326352 308898 326588 309134
rect 332355 309218 332591 309454
rect 332355 308898 332591 309134
rect 430831 309218 431067 309454
rect 430831 308898 431067 309134
rect 434032 309218 434268 309454
rect 434352 309218 434588 309454
rect 434032 308898 434268 309134
rect 434352 308898 434588 309134
rect 448311 309218 448547 309454
rect 448311 308898 448547 309134
rect 546787 309218 547023 309454
rect 546787 308898 547023 309134
rect 571532 309218 571768 309454
rect 571852 309218 572088 309454
rect 571532 308898 571768 309134
rect 571852 308898 572088 309134
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect 9116 291218 9352 291454
rect 9436 291218 9672 291454
rect 9116 290898 9352 291134
rect 9436 290898 9672 291134
rect 56652 291218 56888 291454
rect 56972 291218 57208 291454
rect 56652 290898 56888 291134
rect 56972 290898 57208 291134
rect 92652 291218 92888 291454
rect 92972 291218 93208 291454
rect 92652 290898 92888 291134
rect 92972 290898 93208 291134
rect 128652 291218 128888 291454
rect 128972 291218 129208 291454
rect 128652 290898 128888 291134
rect 128972 290898 129208 291134
rect 164652 291218 164888 291454
rect 164972 291218 165208 291454
rect 164652 290898 164888 291134
rect 164972 290898 165208 291134
rect 200652 291218 200888 291454
rect 200972 291218 201208 291454
rect 200652 290898 200888 291134
rect 200972 290898 201208 291134
rect 236652 291218 236888 291454
rect 236972 291218 237208 291454
rect 236652 290898 236888 291134
rect 236972 290898 237208 291134
rect 272652 291218 272888 291454
rect 272972 291218 273208 291454
rect 272652 290898 272888 291134
rect 272972 290898 273208 291134
rect 308652 291218 308888 291454
rect 308972 291218 309208 291454
rect 308652 290898 308888 291134
rect 308972 290898 309208 291134
rect 344652 291218 344888 291454
rect 344972 291218 345208 291454
rect 344652 290898 344888 291134
rect 344972 290898 345208 291134
rect 380652 291218 380888 291454
rect 380972 291218 381208 291454
rect 380652 290898 380888 291134
rect 380972 290898 381208 291134
rect 416652 291218 416888 291454
rect 416972 291218 417208 291454
rect 416652 290898 416888 291134
rect 416972 290898 417208 291134
rect 452652 291218 452888 291454
rect 452972 291218 453208 291454
rect 452652 290898 452888 291134
rect 452972 290898 453208 291134
rect 488652 291218 488888 291454
rect 488972 291218 489208 291454
rect 488652 290898 488888 291134
rect 488972 290898 489208 291134
rect 524652 291218 524888 291454
rect 524972 291218 525208 291454
rect 524652 290898 524888 291134
rect 524972 290898 525208 291134
rect 560652 291218 560888 291454
rect 560972 291218 561208 291454
rect 560652 290898 560888 291134
rect 560972 290898 561208 291134
rect 570292 291218 570528 291454
rect 570612 291218 570848 291454
rect 570292 290898 570528 291134
rect 570612 290898 570848 291134
rect 7876 273218 8112 273454
rect 8196 273218 8432 273454
rect 7876 272898 8112 273134
rect 8196 272898 8432 273134
rect 38032 273218 38268 273454
rect 38352 273218 38588 273454
rect 38032 272898 38268 273134
rect 38352 272898 38588 273134
rect 74032 273218 74268 273454
rect 74352 273218 74588 273454
rect 74032 272898 74268 273134
rect 74352 272898 74588 273134
rect 110032 273218 110268 273454
rect 110352 273218 110588 273454
rect 110032 272898 110268 273134
rect 110352 272898 110588 273134
rect 146032 273218 146268 273454
rect 146352 273218 146588 273454
rect 146032 272898 146268 273134
rect 146352 272898 146588 273134
rect 182032 273218 182268 273454
rect 182352 273218 182588 273454
rect 182032 272898 182268 273134
rect 182352 272898 182588 273134
rect 218032 273218 218268 273454
rect 218352 273218 218588 273454
rect 218032 272898 218268 273134
rect 218352 272898 218588 273134
rect 254032 273218 254268 273454
rect 254352 273218 254588 273454
rect 254032 272898 254268 273134
rect 254352 272898 254588 273134
rect 290032 273218 290268 273454
rect 290352 273218 290588 273454
rect 290032 272898 290268 273134
rect 290352 272898 290588 273134
rect 326032 273218 326268 273454
rect 326352 273218 326588 273454
rect 326032 272898 326268 273134
rect 326352 272898 326588 273134
rect 362032 273218 362268 273454
rect 362352 273218 362588 273454
rect 362032 272898 362268 273134
rect 362352 272898 362588 273134
rect 398032 273218 398268 273454
rect 398352 273218 398588 273454
rect 398032 272898 398268 273134
rect 398352 272898 398588 273134
rect 434032 273218 434268 273454
rect 434352 273218 434588 273454
rect 434032 272898 434268 273134
rect 434352 272898 434588 273134
rect 470032 273218 470268 273454
rect 470352 273218 470588 273454
rect 470032 272898 470268 273134
rect 470352 272898 470588 273134
rect 506032 273218 506268 273454
rect 506352 273218 506588 273454
rect 506032 272898 506268 273134
rect 506352 272898 506588 273134
rect 542032 273218 542268 273454
rect 542352 273218 542588 273454
rect 542032 272898 542268 273134
rect 542352 272898 542588 273134
rect 571532 273218 571768 273454
rect 571852 273218 572088 273454
rect 571532 272898 571768 273134
rect 571852 272898 572088 273134
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect 9116 255218 9352 255454
rect 9436 255218 9672 255454
rect 9116 254898 9352 255134
rect 9436 254898 9672 255134
rect 56652 255218 56888 255454
rect 56972 255218 57208 255454
rect 56652 254898 56888 255134
rect 56972 254898 57208 255134
rect 92652 255218 92888 255454
rect 92972 255218 93208 255454
rect 92652 254898 92888 255134
rect 92972 254898 93208 255134
rect 128652 255218 128888 255454
rect 128972 255218 129208 255454
rect 128652 254898 128888 255134
rect 128972 254898 129208 255134
rect 164652 255218 164888 255454
rect 164972 255218 165208 255454
rect 164652 254898 164888 255134
rect 164972 254898 165208 255134
rect 200652 255218 200888 255454
rect 200972 255218 201208 255454
rect 200652 254898 200888 255134
rect 200972 254898 201208 255134
rect 236652 255218 236888 255454
rect 236972 255218 237208 255454
rect 236652 254898 236888 255134
rect 236972 254898 237208 255134
rect 272652 255218 272888 255454
rect 272972 255218 273208 255454
rect 272652 254898 272888 255134
rect 272972 254898 273208 255134
rect 308652 255218 308888 255454
rect 308972 255218 309208 255454
rect 308652 254898 308888 255134
rect 308972 254898 309208 255134
rect 344652 255218 344888 255454
rect 344972 255218 345208 255454
rect 344652 254898 344888 255134
rect 344972 254898 345208 255134
rect 380652 255218 380888 255454
rect 380972 255218 381208 255454
rect 380652 254898 380888 255134
rect 380972 254898 381208 255134
rect 416652 255218 416888 255454
rect 416972 255218 417208 255454
rect 416652 254898 416888 255134
rect 416972 254898 417208 255134
rect 452652 255218 452888 255454
rect 452972 255218 453208 255454
rect 452652 254898 452888 255134
rect 452972 254898 453208 255134
rect 488652 255218 488888 255454
rect 488972 255218 489208 255454
rect 488652 254898 488888 255134
rect 488972 254898 489208 255134
rect 524652 255218 524888 255454
rect 524972 255218 525208 255454
rect 524652 254898 524888 255134
rect 524972 254898 525208 255134
rect 560652 255218 560888 255454
rect 560972 255218 561208 255454
rect 560652 254898 560888 255134
rect 560972 254898 561208 255134
rect 570292 255218 570528 255454
rect 570612 255218 570848 255454
rect 570292 254898 570528 255134
rect 570612 254898 570848 255134
rect 7876 237218 8112 237454
rect 8196 237218 8432 237454
rect 7876 236898 8112 237134
rect 8196 236898 8432 237134
rect 38032 237218 38268 237454
rect 38352 237218 38588 237454
rect 38032 236898 38268 237134
rect 38352 236898 38588 237134
rect 74032 237218 74268 237454
rect 74352 237218 74588 237454
rect 74032 236898 74268 237134
rect 74352 236898 74588 237134
rect 110032 237218 110268 237454
rect 110352 237218 110588 237454
rect 110032 236898 110268 237134
rect 110352 236898 110588 237134
rect 146032 237218 146268 237454
rect 146352 237218 146588 237454
rect 146032 236898 146268 237134
rect 146352 236898 146588 237134
rect 182032 237218 182268 237454
rect 182352 237218 182588 237454
rect 182032 236898 182268 237134
rect 182352 236898 182588 237134
rect 218032 237218 218268 237454
rect 218352 237218 218588 237454
rect 218032 236898 218268 237134
rect 218352 236898 218588 237134
rect 254032 237218 254268 237454
rect 254352 237218 254588 237454
rect 254032 236898 254268 237134
rect 254352 236898 254588 237134
rect 290032 237218 290268 237454
rect 290352 237218 290588 237454
rect 290032 236898 290268 237134
rect 290352 236898 290588 237134
rect 326032 237218 326268 237454
rect 326352 237218 326588 237454
rect 326032 236898 326268 237134
rect 326352 236898 326588 237134
rect 362032 237218 362268 237454
rect 362352 237218 362588 237454
rect 362032 236898 362268 237134
rect 362352 236898 362588 237134
rect 398032 237218 398268 237454
rect 398352 237218 398588 237454
rect 398032 236898 398268 237134
rect 398352 236898 398588 237134
rect 434032 237218 434268 237454
rect 434352 237218 434588 237454
rect 434032 236898 434268 237134
rect 434352 236898 434588 237134
rect 470032 237218 470268 237454
rect 470352 237218 470588 237454
rect 470032 236898 470268 237134
rect 470352 236898 470588 237134
rect 506032 237218 506268 237454
rect 506352 237218 506588 237454
rect 506032 236898 506268 237134
rect 506352 236898 506588 237134
rect 542032 237218 542268 237454
rect 542352 237218 542588 237454
rect 542032 236898 542268 237134
rect 542352 236898 542588 237134
rect 571532 237218 571768 237454
rect 571852 237218 572088 237454
rect 571532 236898 571768 237134
rect 571852 236898 572088 237134
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect 9116 219218 9352 219454
rect 9436 219218 9672 219454
rect 9116 218898 9352 219134
rect 9436 218898 9672 219134
rect 56652 219218 56888 219454
rect 56972 219218 57208 219454
rect 56652 218898 56888 219134
rect 56972 218898 57208 219134
rect 92652 219218 92888 219454
rect 92972 219218 93208 219454
rect 92652 218898 92888 219134
rect 92972 218898 93208 219134
rect 128652 219218 128888 219454
rect 128972 219218 129208 219454
rect 128652 218898 128888 219134
rect 128972 218898 129208 219134
rect 164652 219218 164888 219454
rect 164972 219218 165208 219454
rect 164652 218898 164888 219134
rect 164972 218898 165208 219134
rect 200652 219218 200888 219454
rect 200972 219218 201208 219454
rect 200652 218898 200888 219134
rect 200972 218898 201208 219134
rect 236652 219218 236888 219454
rect 236972 219218 237208 219454
rect 236652 218898 236888 219134
rect 236972 218898 237208 219134
rect 272652 219218 272888 219454
rect 272972 219218 273208 219454
rect 272652 218898 272888 219134
rect 272972 218898 273208 219134
rect 308652 219218 308888 219454
rect 308972 219218 309208 219454
rect 308652 218898 308888 219134
rect 308972 218898 309208 219134
rect 344652 219218 344888 219454
rect 344972 219218 345208 219454
rect 344652 218898 344888 219134
rect 344972 218898 345208 219134
rect 380652 219218 380888 219454
rect 380972 219218 381208 219454
rect 380652 218898 380888 219134
rect 380972 218898 381208 219134
rect 416652 219218 416888 219454
rect 416972 219218 417208 219454
rect 416652 218898 416888 219134
rect 416972 218898 417208 219134
rect 452652 219218 452888 219454
rect 452972 219218 453208 219454
rect 452652 218898 452888 219134
rect 452972 218898 453208 219134
rect 488652 219218 488888 219454
rect 488972 219218 489208 219454
rect 488652 218898 488888 219134
rect 488972 218898 489208 219134
rect 524652 219218 524888 219454
rect 524972 219218 525208 219454
rect 524652 218898 524888 219134
rect 524972 218898 525208 219134
rect 560652 219218 560888 219454
rect 560972 219218 561208 219454
rect 560652 218898 560888 219134
rect 560972 218898 561208 219134
rect 570292 219218 570528 219454
rect 570612 219218 570848 219454
rect 570292 218898 570528 219134
rect 570612 218898 570848 219134
rect 7876 201218 8112 201454
rect 8196 201218 8432 201454
rect 7876 200898 8112 201134
rect 8196 200898 8432 201134
rect 38032 201218 38268 201454
rect 38352 201218 38588 201454
rect 38032 200898 38268 201134
rect 38352 200898 38588 201134
rect 74032 201218 74268 201454
rect 74352 201218 74588 201454
rect 74032 200898 74268 201134
rect 74352 200898 74588 201134
rect 110032 201218 110268 201454
rect 110352 201218 110588 201454
rect 110032 200898 110268 201134
rect 110352 200898 110588 201134
rect 146032 201218 146268 201454
rect 146352 201218 146588 201454
rect 146032 200898 146268 201134
rect 146352 200898 146588 201134
rect 182032 201218 182268 201454
rect 182352 201218 182588 201454
rect 182032 200898 182268 201134
rect 182352 200898 182588 201134
rect 218032 201218 218268 201454
rect 218352 201218 218588 201454
rect 218032 200898 218268 201134
rect 218352 200898 218588 201134
rect 254032 201218 254268 201454
rect 254352 201218 254588 201454
rect 254032 200898 254268 201134
rect 254352 200898 254588 201134
rect 290032 201218 290268 201454
rect 290352 201218 290588 201454
rect 290032 200898 290268 201134
rect 290352 200898 290588 201134
rect 326032 201218 326268 201454
rect 326352 201218 326588 201454
rect 326032 200898 326268 201134
rect 326352 200898 326588 201134
rect 362032 201218 362268 201454
rect 362352 201218 362588 201454
rect 362032 200898 362268 201134
rect 362352 200898 362588 201134
rect 398032 201218 398268 201454
rect 398352 201218 398588 201454
rect 398032 200898 398268 201134
rect 398352 200898 398588 201134
rect 434032 201218 434268 201454
rect 434352 201218 434588 201454
rect 434032 200898 434268 201134
rect 434352 200898 434588 201134
rect 470032 201218 470268 201454
rect 470352 201218 470588 201454
rect 470032 200898 470268 201134
rect 470352 200898 470588 201134
rect 506032 201218 506268 201454
rect 506352 201218 506588 201454
rect 506032 200898 506268 201134
rect 506352 200898 506588 201134
rect 542032 201218 542268 201454
rect 542352 201218 542588 201454
rect 542032 200898 542268 201134
rect 542352 200898 542588 201134
rect 571532 201218 571768 201454
rect 571852 201218 572088 201454
rect 571532 200898 571768 201134
rect 571852 200898 572088 201134
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect 9116 183218 9352 183454
rect 9436 183218 9672 183454
rect 9116 182898 9352 183134
rect 9436 182898 9672 183134
rect 56652 183218 56888 183454
rect 56972 183218 57208 183454
rect 56652 182898 56888 183134
rect 56972 182898 57208 183134
rect 92652 183218 92888 183454
rect 92972 183218 93208 183454
rect 92652 182898 92888 183134
rect 92972 182898 93208 183134
rect 128652 183218 128888 183454
rect 128972 183218 129208 183454
rect 128652 182898 128888 183134
rect 128972 182898 129208 183134
rect 164652 183218 164888 183454
rect 164972 183218 165208 183454
rect 164652 182898 164888 183134
rect 164972 182898 165208 183134
rect 200652 183218 200888 183454
rect 200972 183218 201208 183454
rect 200652 182898 200888 183134
rect 200972 182898 201208 183134
rect 236652 183218 236888 183454
rect 236972 183218 237208 183454
rect 236652 182898 236888 183134
rect 236972 182898 237208 183134
rect 272652 183218 272888 183454
rect 272972 183218 273208 183454
rect 272652 182898 272888 183134
rect 272972 182898 273208 183134
rect 308652 183218 308888 183454
rect 308972 183218 309208 183454
rect 308652 182898 308888 183134
rect 308972 182898 309208 183134
rect 344652 183218 344888 183454
rect 344972 183218 345208 183454
rect 344652 182898 344888 183134
rect 344972 182898 345208 183134
rect 380652 183218 380888 183454
rect 380972 183218 381208 183454
rect 380652 182898 380888 183134
rect 380972 182898 381208 183134
rect 416652 183218 416888 183454
rect 416972 183218 417208 183454
rect 416652 182898 416888 183134
rect 416972 182898 417208 183134
rect 452652 183218 452888 183454
rect 452972 183218 453208 183454
rect 452652 182898 452888 183134
rect 452972 182898 453208 183134
rect 488652 183218 488888 183454
rect 488972 183218 489208 183454
rect 488652 182898 488888 183134
rect 488972 182898 489208 183134
rect 524652 183218 524888 183454
rect 524972 183218 525208 183454
rect 524652 182898 524888 183134
rect 524972 182898 525208 183134
rect 560652 183218 560888 183454
rect 560972 183218 561208 183454
rect 560652 182898 560888 183134
rect 560972 182898 561208 183134
rect 570292 183218 570528 183454
rect 570612 183218 570848 183454
rect 570292 182898 570528 183134
rect 570612 182898 570848 183134
rect 7876 165218 8112 165454
rect 8196 165218 8432 165454
rect 7876 164898 8112 165134
rect 8196 164898 8432 165134
rect 38032 165218 38268 165454
rect 38352 165218 38588 165454
rect 38032 164898 38268 165134
rect 38352 164898 38588 165134
rect 74032 165218 74268 165454
rect 74352 165218 74588 165454
rect 74032 164898 74268 165134
rect 74352 164898 74588 165134
rect 110032 165218 110268 165454
rect 110352 165218 110588 165454
rect 110032 164898 110268 165134
rect 110352 164898 110588 165134
rect 146032 165218 146268 165454
rect 146352 165218 146588 165454
rect 146032 164898 146268 165134
rect 146352 164898 146588 165134
rect 182032 165218 182268 165454
rect 182352 165218 182588 165454
rect 182032 164898 182268 165134
rect 182352 164898 182588 165134
rect 218032 165218 218268 165454
rect 218352 165218 218588 165454
rect 218032 164898 218268 165134
rect 218352 164898 218588 165134
rect 254032 165218 254268 165454
rect 254352 165218 254588 165454
rect 254032 164898 254268 165134
rect 254352 164898 254588 165134
rect 290032 165218 290268 165454
rect 290352 165218 290588 165454
rect 290032 164898 290268 165134
rect 290352 164898 290588 165134
rect 326032 165218 326268 165454
rect 326352 165218 326588 165454
rect 326032 164898 326268 165134
rect 326352 164898 326588 165134
rect 362032 165218 362268 165454
rect 362352 165218 362588 165454
rect 362032 164898 362268 165134
rect 362352 164898 362588 165134
rect 398032 165218 398268 165454
rect 398352 165218 398588 165454
rect 398032 164898 398268 165134
rect 398352 164898 398588 165134
rect 434032 165218 434268 165454
rect 434352 165218 434588 165454
rect 434032 164898 434268 165134
rect 434352 164898 434588 165134
rect 470032 165218 470268 165454
rect 470352 165218 470588 165454
rect 470032 164898 470268 165134
rect 470352 164898 470588 165134
rect 506032 165218 506268 165454
rect 506352 165218 506588 165454
rect 506032 164898 506268 165134
rect 506352 164898 506588 165134
rect 542032 165218 542268 165454
rect 542352 165218 542588 165454
rect 542032 164898 542268 165134
rect 542352 164898 542588 165134
rect 571532 165218 571768 165454
rect 571852 165218 572088 165454
rect 571532 164898 571768 165134
rect 571852 164898 572088 165134
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect 9116 147218 9352 147454
rect 9436 147218 9672 147454
rect 9116 146898 9352 147134
rect 9436 146898 9672 147134
rect 56652 147218 56888 147454
rect 56972 147218 57208 147454
rect 56652 146898 56888 147134
rect 56972 146898 57208 147134
rect 92652 147218 92888 147454
rect 92972 147218 93208 147454
rect 92652 146898 92888 147134
rect 92972 146898 93208 147134
rect 128652 147218 128888 147454
rect 128972 147218 129208 147454
rect 128652 146898 128888 147134
rect 128972 146898 129208 147134
rect 164652 147218 164888 147454
rect 164972 147218 165208 147454
rect 164652 146898 164888 147134
rect 164972 146898 165208 147134
rect 200652 147218 200888 147454
rect 200972 147218 201208 147454
rect 200652 146898 200888 147134
rect 200972 146898 201208 147134
rect 236652 147218 236888 147454
rect 236972 147218 237208 147454
rect 236652 146898 236888 147134
rect 236972 146898 237208 147134
rect 272652 147218 272888 147454
rect 272972 147218 273208 147454
rect 272652 146898 272888 147134
rect 272972 146898 273208 147134
rect 308652 147218 308888 147454
rect 308972 147218 309208 147454
rect 308652 146898 308888 147134
rect 308972 146898 309208 147134
rect 344652 147218 344888 147454
rect 344972 147218 345208 147454
rect 344652 146898 344888 147134
rect 344972 146898 345208 147134
rect 380652 147218 380888 147454
rect 380972 147218 381208 147454
rect 380652 146898 380888 147134
rect 380972 146898 381208 147134
rect 416652 147218 416888 147454
rect 416972 147218 417208 147454
rect 416652 146898 416888 147134
rect 416972 146898 417208 147134
rect 452652 147218 452888 147454
rect 452972 147218 453208 147454
rect 452652 146898 452888 147134
rect 452972 146898 453208 147134
rect 488652 147218 488888 147454
rect 488972 147218 489208 147454
rect 488652 146898 488888 147134
rect 488972 146898 489208 147134
rect 524652 147218 524888 147454
rect 524972 147218 525208 147454
rect 524652 146898 524888 147134
rect 524972 146898 525208 147134
rect 560652 147218 560888 147454
rect 560972 147218 561208 147454
rect 560652 146898 560888 147134
rect 560972 146898 561208 147134
rect 570292 147218 570528 147454
rect 570612 147218 570848 147454
rect 570292 146898 570528 147134
rect 570612 146898 570848 147134
rect 7876 129218 8112 129454
rect 8196 129218 8432 129454
rect 7876 128898 8112 129134
rect 8196 128898 8432 129134
rect 38032 129218 38268 129454
rect 38352 129218 38588 129454
rect 38032 128898 38268 129134
rect 38352 128898 38588 129134
rect 74032 129218 74268 129454
rect 74352 129218 74588 129454
rect 74032 128898 74268 129134
rect 74352 128898 74588 129134
rect 110032 129218 110268 129454
rect 110352 129218 110588 129454
rect 110032 128898 110268 129134
rect 110352 128898 110588 129134
rect 146032 129218 146268 129454
rect 146352 129218 146588 129454
rect 146032 128898 146268 129134
rect 146352 128898 146588 129134
rect 182032 129218 182268 129454
rect 182352 129218 182588 129454
rect 182032 128898 182268 129134
rect 182352 128898 182588 129134
rect 218032 129218 218268 129454
rect 218352 129218 218588 129454
rect 218032 128898 218268 129134
rect 218352 128898 218588 129134
rect 254032 129218 254268 129454
rect 254352 129218 254588 129454
rect 254032 128898 254268 129134
rect 254352 128898 254588 129134
rect 290032 129218 290268 129454
rect 290352 129218 290588 129454
rect 290032 128898 290268 129134
rect 290352 128898 290588 129134
rect 326032 129218 326268 129454
rect 326352 129218 326588 129454
rect 326032 128898 326268 129134
rect 326352 128898 326588 129134
rect 362032 129218 362268 129454
rect 362352 129218 362588 129454
rect 362032 128898 362268 129134
rect 362352 128898 362588 129134
rect 398032 129218 398268 129454
rect 398352 129218 398588 129454
rect 398032 128898 398268 129134
rect 398352 128898 398588 129134
rect 434032 129218 434268 129454
rect 434352 129218 434588 129454
rect 434032 128898 434268 129134
rect 434352 128898 434588 129134
rect 470032 129218 470268 129454
rect 470352 129218 470588 129454
rect 470032 128898 470268 129134
rect 470352 128898 470588 129134
rect 506032 129218 506268 129454
rect 506352 129218 506588 129454
rect 506032 128898 506268 129134
rect 506352 128898 506588 129134
rect 542032 129218 542268 129454
rect 542352 129218 542588 129454
rect 542032 128898 542268 129134
rect 542352 128898 542588 129134
rect 571532 129218 571768 129454
rect 571852 129218 572088 129454
rect 571532 128898 571768 129134
rect 571852 128898 572088 129134
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect 9116 111218 9352 111454
rect 9436 111218 9672 111454
rect 9116 110898 9352 111134
rect 9436 110898 9672 111134
rect 56652 111218 56888 111454
rect 56972 111218 57208 111454
rect 56652 110898 56888 111134
rect 56972 110898 57208 111134
rect 92652 111218 92888 111454
rect 92972 111218 93208 111454
rect 92652 110898 92888 111134
rect 92972 110898 93208 111134
rect 128652 111218 128888 111454
rect 128972 111218 129208 111454
rect 128652 110898 128888 111134
rect 128972 110898 129208 111134
rect 164652 111218 164888 111454
rect 164972 111218 165208 111454
rect 164652 110898 164888 111134
rect 164972 110898 165208 111134
rect 200652 111218 200888 111454
rect 200972 111218 201208 111454
rect 200652 110898 200888 111134
rect 200972 110898 201208 111134
rect 236652 111218 236888 111454
rect 236972 111218 237208 111454
rect 236652 110898 236888 111134
rect 236972 110898 237208 111134
rect 272652 111218 272888 111454
rect 272972 111218 273208 111454
rect 272652 110898 272888 111134
rect 272972 110898 273208 111134
rect 308652 111218 308888 111454
rect 308972 111218 309208 111454
rect 308652 110898 308888 111134
rect 308972 110898 309208 111134
rect 344652 111218 344888 111454
rect 344972 111218 345208 111454
rect 344652 110898 344888 111134
rect 344972 110898 345208 111134
rect 380652 111218 380888 111454
rect 380972 111218 381208 111454
rect 380652 110898 380888 111134
rect 380972 110898 381208 111134
rect 416652 111218 416888 111454
rect 416972 111218 417208 111454
rect 416652 110898 416888 111134
rect 416972 110898 417208 111134
rect 452652 111218 452888 111454
rect 452972 111218 453208 111454
rect 452652 110898 452888 111134
rect 452972 110898 453208 111134
rect 488652 111218 488888 111454
rect 488972 111218 489208 111454
rect 488652 110898 488888 111134
rect 488972 110898 489208 111134
rect 524652 111218 524888 111454
rect 524972 111218 525208 111454
rect 524652 110898 524888 111134
rect 524972 110898 525208 111134
rect 560652 111218 560888 111454
rect 560972 111218 561208 111454
rect 560652 110898 560888 111134
rect 560972 110898 561208 111134
rect 570292 111218 570528 111454
rect 570612 111218 570848 111454
rect 570292 110898 570528 111134
rect 570612 110898 570848 111134
rect 7876 93218 8112 93454
rect 8196 93218 8432 93454
rect 7876 92898 8112 93134
rect 8196 92898 8432 93134
rect 38032 93218 38268 93454
rect 38352 93218 38588 93454
rect 38032 92898 38268 93134
rect 38352 92898 38588 93134
rect 74032 93218 74268 93454
rect 74352 93218 74588 93454
rect 74032 92898 74268 93134
rect 74352 92898 74588 93134
rect 110032 93218 110268 93454
rect 110352 93218 110588 93454
rect 110032 92898 110268 93134
rect 110352 92898 110588 93134
rect 146032 93218 146268 93454
rect 146352 93218 146588 93454
rect 146032 92898 146268 93134
rect 146352 92898 146588 93134
rect 182032 93218 182268 93454
rect 182352 93218 182588 93454
rect 182032 92898 182268 93134
rect 182352 92898 182588 93134
rect 218032 93218 218268 93454
rect 218352 93218 218588 93454
rect 218032 92898 218268 93134
rect 218352 92898 218588 93134
rect 254032 93218 254268 93454
rect 254352 93218 254588 93454
rect 254032 92898 254268 93134
rect 254352 92898 254588 93134
rect 290032 93218 290268 93454
rect 290352 93218 290588 93454
rect 290032 92898 290268 93134
rect 290352 92898 290588 93134
rect 326032 93218 326268 93454
rect 326352 93218 326588 93454
rect 326032 92898 326268 93134
rect 326352 92898 326588 93134
rect 362032 93218 362268 93454
rect 362352 93218 362588 93454
rect 362032 92898 362268 93134
rect 362352 92898 362588 93134
rect 398032 93218 398268 93454
rect 398352 93218 398588 93454
rect 398032 92898 398268 93134
rect 398352 92898 398588 93134
rect 434032 93218 434268 93454
rect 434352 93218 434588 93454
rect 434032 92898 434268 93134
rect 434352 92898 434588 93134
rect 470032 93218 470268 93454
rect 470352 93218 470588 93454
rect 470032 92898 470268 93134
rect 470352 92898 470588 93134
rect 506032 93218 506268 93454
rect 506352 93218 506588 93454
rect 506032 92898 506268 93134
rect 506352 92898 506588 93134
rect 542032 93218 542268 93454
rect 542352 93218 542588 93454
rect 542032 92898 542268 93134
rect 542352 92898 542588 93134
rect 571532 93218 571768 93454
rect 571852 93218 572088 93454
rect 571532 92898 571768 93134
rect 571852 92898 572088 93134
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect 9116 75218 9352 75454
rect 9436 75218 9672 75454
rect 9116 74898 9352 75134
rect 9436 74898 9672 75134
rect 56652 75218 56888 75454
rect 56972 75218 57208 75454
rect 56652 74898 56888 75134
rect 56972 74898 57208 75134
rect 92652 75218 92888 75454
rect 92972 75218 93208 75454
rect 92652 74898 92888 75134
rect 92972 74898 93208 75134
rect 128652 75218 128888 75454
rect 128972 75218 129208 75454
rect 128652 74898 128888 75134
rect 128972 74898 129208 75134
rect 164652 75218 164888 75454
rect 164972 75218 165208 75454
rect 164652 74898 164888 75134
rect 164972 74898 165208 75134
rect 200652 75218 200888 75454
rect 200972 75218 201208 75454
rect 200652 74898 200888 75134
rect 200972 74898 201208 75134
rect 236652 75218 236888 75454
rect 236972 75218 237208 75454
rect 236652 74898 236888 75134
rect 236972 74898 237208 75134
rect 272652 75218 272888 75454
rect 272972 75218 273208 75454
rect 272652 74898 272888 75134
rect 272972 74898 273208 75134
rect 308652 75218 308888 75454
rect 308972 75218 309208 75454
rect 308652 74898 308888 75134
rect 308972 74898 309208 75134
rect 344652 75218 344888 75454
rect 344972 75218 345208 75454
rect 344652 74898 344888 75134
rect 344972 74898 345208 75134
rect 380652 75218 380888 75454
rect 380972 75218 381208 75454
rect 380652 74898 380888 75134
rect 380972 74898 381208 75134
rect 416652 75218 416888 75454
rect 416972 75218 417208 75454
rect 416652 74898 416888 75134
rect 416972 74898 417208 75134
rect 452652 75218 452888 75454
rect 452972 75218 453208 75454
rect 452652 74898 452888 75134
rect 452972 74898 453208 75134
rect 488652 75218 488888 75454
rect 488972 75218 489208 75454
rect 488652 74898 488888 75134
rect 488972 74898 489208 75134
rect 524652 75218 524888 75454
rect 524972 75218 525208 75454
rect 524652 74898 524888 75134
rect 524972 74898 525208 75134
rect 560652 75218 560888 75454
rect 560972 75218 561208 75454
rect 560652 74898 560888 75134
rect 560972 74898 561208 75134
rect 570292 75218 570528 75454
rect 570612 75218 570848 75454
rect 570292 74898 570528 75134
rect 570612 74898 570848 75134
rect 7876 57218 8112 57454
rect 8196 57218 8432 57454
rect 7876 56898 8112 57134
rect 8196 56898 8432 57134
rect 38032 57218 38268 57454
rect 38352 57218 38588 57454
rect 38032 56898 38268 57134
rect 38352 56898 38588 57134
rect 74032 57218 74268 57454
rect 74352 57218 74588 57454
rect 74032 56898 74268 57134
rect 74352 56898 74588 57134
rect 110032 57218 110268 57454
rect 110352 57218 110588 57454
rect 110032 56898 110268 57134
rect 110352 56898 110588 57134
rect 146032 57218 146268 57454
rect 146352 57218 146588 57454
rect 146032 56898 146268 57134
rect 146352 56898 146588 57134
rect 182032 57218 182268 57454
rect 182352 57218 182588 57454
rect 182032 56898 182268 57134
rect 182352 56898 182588 57134
rect 218032 57218 218268 57454
rect 218352 57218 218588 57454
rect 218032 56898 218268 57134
rect 218352 56898 218588 57134
rect 254032 57218 254268 57454
rect 254352 57218 254588 57454
rect 254032 56898 254268 57134
rect 254352 56898 254588 57134
rect 290032 57218 290268 57454
rect 290352 57218 290588 57454
rect 290032 56898 290268 57134
rect 290352 56898 290588 57134
rect 326032 57218 326268 57454
rect 326352 57218 326588 57454
rect 326032 56898 326268 57134
rect 326352 56898 326588 57134
rect 362032 57218 362268 57454
rect 362352 57218 362588 57454
rect 362032 56898 362268 57134
rect 362352 56898 362588 57134
rect 398032 57218 398268 57454
rect 398352 57218 398588 57454
rect 398032 56898 398268 57134
rect 398352 56898 398588 57134
rect 434032 57218 434268 57454
rect 434352 57218 434588 57454
rect 434032 56898 434268 57134
rect 434352 56898 434588 57134
rect 470032 57218 470268 57454
rect 470352 57218 470588 57454
rect 470032 56898 470268 57134
rect 470352 56898 470588 57134
rect 506032 57218 506268 57454
rect 506352 57218 506588 57454
rect 506032 56898 506268 57134
rect 506352 56898 506588 57134
rect 542032 57218 542268 57454
rect 542352 57218 542588 57454
rect 542032 56898 542268 57134
rect 542352 56898 542588 57134
rect 571532 57218 571768 57454
rect 571852 57218 572088 57454
rect 571532 56898 571768 57134
rect 571852 56898 572088 57134
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect 9116 39218 9352 39454
rect 9436 39218 9672 39454
rect 9116 38898 9352 39134
rect 9436 38898 9672 39134
rect 56652 39218 56888 39454
rect 56972 39218 57208 39454
rect 56652 38898 56888 39134
rect 56972 38898 57208 39134
rect 92652 39218 92888 39454
rect 92972 39218 93208 39454
rect 92652 38898 92888 39134
rect 92972 38898 93208 39134
rect 128652 39218 128888 39454
rect 128972 39218 129208 39454
rect 128652 38898 128888 39134
rect 128972 38898 129208 39134
rect 164652 39218 164888 39454
rect 164972 39218 165208 39454
rect 164652 38898 164888 39134
rect 164972 38898 165208 39134
rect 200652 39218 200888 39454
rect 200972 39218 201208 39454
rect 200652 38898 200888 39134
rect 200972 38898 201208 39134
rect 236652 39218 236888 39454
rect 236972 39218 237208 39454
rect 236652 38898 236888 39134
rect 236972 38898 237208 39134
rect 272652 39218 272888 39454
rect 272972 39218 273208 39454
rect 272652 38898 272888 39134
rect 272972 38898 273208 39134
rect 308652 39218 308888 39454
rect 308972 39218 309208 39454
rect 308652 38898 308888 39134
rect 308972 38898 309208 39134
rect 344652 39218 344888 39454
rect 344972 39218 345208 39454
rect 344652 38898 344888 39134
rect 344972 38898 345208 39134
rect 380652 39218 380888 39454
rect 380972 39218 381208 39454
rect 380652 38898 380888 39134
rect 380972 38898 381208 39134
rect 416652 39218 416888 39454
rect 416972 39218 417208 39454
rect 416652 38898 416888 39134
rect 416972 38898 417208 39134
rect 452652 39218 452888 39454
rect 452972 39218 453208 39454
rect 452652 38898 452888 39134
rect 452972 38898 453208 39134
rect 488652 39218 488888 39454
rect 488972 39218 489208 39454
rect 488652 38898 488888 39134
rect 488972 38898 489208 39134
rect 524652 39218 524888 39454
rect 524972 39218 525208 39454
rect 524652 38898 524888 39134
rect 524972 38898 525208 39134
rect 560652 39218 560888 39454
rect 560972 39218 561208 39454
rect 560652 38898 560888 39134
rect 560972 38898 561208 39134
rect 570292 39218 570528 39454
rect 570612 39218 570848 39454
rect 570292 38898 570528 39134
rect 570612 38898 570848 39134
rect 7876 21218 8112 21454
rect 8196 21218 8432 21454
rect 7876 20898 8112 21134
rect 8196 20898 8432 21134
rect 38032 21218 38268 21454
rect 38352 21218 38588 21454
rect 38032 20898 38268 21134
rect 38352 20898 38588 21134
rect 74032 21218 74268 21454
rect 74352 21218 74588 21454
rect 74032 20898 74268 21134
rect 74352 20898 74588 21134
rect 110032 21218 110268 21454
rect 110352 21218 110588 21454
rect 110032 20898 110268 21134
rect 110352 20898 110588 21134
rect 146032 21218 146268 21454
rect 146352 21218 146588 21454
rect 146032 20898 146268 21134
rect 146352 20898 146588 21134
rect 182032 21218 182268 21454
rect 182352 21218 182588 21454
rect 182032 20898 182268 21134
rect 182352 20898 182588 21134
rect 218032 21218 218268 21454
rect 218352 21218 218588 21454
rect 218032 20898 218268 21134
rect 218352 20898 218588 21134
rect 254032 21218 254268 21454
rect 254352 21218 254588 21454
rect 254032 20898 254268 21134
rect 254352 20898 254588 21134
rect 290032 21218 290268 21454
rect 290352 21218 290588 21454
rect 290032 20898 290268 21134
rect 290352 20898 290588 21134
rect 326032 21218 326268 21454
rect 326352 21218 326588 21454
rect 326032 20898 326268 21134
rect 326352 20898 326588 21134
rect 362032 21218 362268 21454
rect 362352 21218 362588 21454
rect 362032 20898 362268 21134
rect 362352 20898 362588 21134
rect 398032 21218 398268 21454
rect 398352 21218 398588 21454
rect 398032 20898 398268 21134
rect 398352 20898 398588 21134
rect 434032 21218 434268 21454
rect 434352 21218 434588 21454
rect 434032 20898 434268 21134
rect 434352 20898 434588 21134
rect 470032 21218 470268 21454
rect 470352 21218 470588 21454
rect 470032 20898 470268 21134
rect 470352 20898 470588 21134
rect 506032 21218 506268 21454
rect 506352 21218 506588 21454
rect 506032 20898 506268 21134
rect 506352 20898 506588 21134
rect 542032 21218 542268 21454
rect 542352 21218 542588 21454
rect 542032 20898 542268 21134
rect 542352 20898 542588 21134
rect 571532 21218 571768 21454
rect 571852 21218 572088 21454
rect 571532 20898 571768 21134
rect 571852 20898 572088 21134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 9116 687454
rect 9352 687218 9436 687454
rect 9672 687218 56652 687454
rect 56888 687218 56972 687454
rect 57208 687218 92652 687454
rect 92888 687218 92972 687454
rect 93208 687218 128652 687454
rect 128888 687218 128972 687454
rect 129208 687218 164652 687454
rect 164888 687218 164972 687454
rect 165208 687218 200652 687454
rect 200888 687218 200972 687454
rect 201208 687218 236652 687454
rect 236888 687218 236972 687454
rect 237208 687218 272652 687454
rect 272888 687218 272972 687454
rect 273208 687218 308652 687454
rect 308888 687218 308972 687454
rect 309208 687218 344652 687454
rect 344888 687218 344972 687454
rect 345208 687218 380652 687454
rect 380888 687218 380972 687454
rect 381208 687218 416652 687454
rect 416888 687218 416972 687454
rect 417208 687218 452652 687454
rect 452888 687218 452972 687454
rect 453208 687218 488652 687454
rect 488888 687218 488972 687454
rect 489208 687218 524652 687454
rect 524888 687218 524972 687454
rect 525208 687218 560652 687454
rect 560888 687218 560972 687454
rect 561208 687218 570292 687454
rect 570528 687218 570612 687454
rect 570848 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 9116 687134
rect 9352 686898 9436 687134
rect 9672 686898 56652 687134
rect 56888 686898 56972 687134
rect 57208 686898 92652 687134
rect 92888 686898 92972 687134
rect 93208 686898 128652 687134
rect 128888 686898 128972 687134
rect 129208 686898 164652 687134
rect 164888 686898 164972 687134
rect 165208 686898 200652 687134
rect 200888 686898 200972 687134
rect 201208 686898 236652 687134
rect 236888 686898 236972 687134
rect 237208 686898 272652 687134
rect 272888 686898 272972 687134
rect 273208 686898 308652 687134
rect 308888 686898 308972 687134
rect 309208 686898 344652 687134
rect 344888 686898 344972 687134
rect 345208 686898 380652 687134
rect 380888 686898 380972 687134
rect 381208 686898 416652 687134
rect 416888 686898 416972 687134
rect 417208 686898 452652 687134
rect 452888 686898 452972 687134
rect 453208 686898 488652 687134
rect 488888 686898 488972 687134
rect 489208 686898 524652 687134
rect 524888 686898 524972 687134
rect 525208 686898 560652 687134
rect 560888 686898 560972 687134
rect 561208 686898 570292 687134
rect 570528 686898 570612 687134
rect 570848 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 7876 669454
rect 8112 669218 8196 669454
rect 8432 669218 38032 669454
rect 38268 669218 38352 669454
rect 38588 669218 74032 669454
rect 74268 669218 74352 669454
rect 74588 669218 100443 669454
rect 100679 669218 198919 669454
rect 199155 669218 216399 669454
rect 216635 669218 314875 669454
rect 315111 669218 326032 669454
rect 326268 669218 326352 669454
rect 326588 669218 332355 669454
rect 332591 669218 430831 669454
rect 431067 669218 434032 669454
rect 434268 669218 434352 669454
rect 434588 669218 448311 669454
rect 448547 669218 546787 669454
rect 547023 669218 571532 669454
rect 571768 669218 571852 669454
rect 572088 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 7876 669134
rect 8112 668898 8196 669134
rect 8432 668898 38032 669134
rect 38268 668898 38352 669134
rect 38588 668898 74032 669134
rect 74268 668898 74352 669134
rect 74588 668898 100443 669134
rect 100679 668898 198919 669134
rect 199155 668898 216399 669134
rect 216635 668898 314875 669134
rect 315111 668898 326032 669134
rect 326268 668898 326352 669134
rect 326588 668898 332355 669134
rect 332591 668898 430831 669134
rect 431067 668898 434032 669134
rect 434268 668898 434352 669134
rect 434588 668898 448311 669134
rect 448547 668898 546787 669134
rect 547023 668898 571532 669134
rect 571768 668898 571852 669134
rect 572088 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 9116 651454
rect 9352 651218 9436 651454
rect 9672 651218 56652 651454
rect 56888 651218 56972 651454
rect 57208 651218 92652 651454
rect 92888 651218 92972 651454
rect 93208 651218 101163 651454
rect 101399 651218 198199 651454
rect 198435 651218 200652 651454
rect 200888 651218 200972 651454
rect 201208 651218 217119 651454
rect 217355 651218 314155 651454
rect 314391 651218 333075 651454
rect 333311 651218 430111 651454
rect 430347 651218 449031 651454
rect 449267 651218 546067 651454
rect 546303 651218 560652 651454
rect 560888 651218 560972 651454
rect 561208 651218 570292 651454
rect 570528 651218 570612 651454
rect 570848 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 9116 651134
rect 9352 650898 9436 651134
rect 9672 650898 56652 651134
rect 56888 650898 56972 651134
rect 57208 650898 92652 651134
rect 92888 650898 92972 651134
rect 93208 650898 101163 651134
rect 101399 650898 198199 651134
rect 198435 650898 200652 651134
rect 200888 650898 200972 651134
rect 201208 650898 217119 651134
rect 217355 650898 314155 651134
rect 314391 650898 333075 651134
rect 333311 650898 430111 651134
rect 430347 650898 449031 651134
rect 449267 650898 546067 651134
rect 546303 650898 560652 651134
rect 560888 650898 560972 651134
rect 561208 650898 570292 651134
rect 570528 650898 570612 651134
rect 570848 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 7876 633454
rect 8112 633218 8196 633454
rect 8432 633218 38032 633454
rect 38268 633218 38352 633454
rect 38588 633218 74032 633454
rect 74268 633218 74352 633454
rect 74588 633218 100443 633454
rect 100679 633218 198919 633454
rect 199155 633218 216399 633454
rect 216635 633218 314875 633454
rect 315111 633218 326032 633454
rect 326268 633218 326352 633454
rect 326588 633218 332355 633454
rect 332591 633218 430831 633454
rect 431067 633218 434032 633454
rect 434268 633218 434352 633454
rect 434588 633218 448311 633454
rect 448547 633218 546787 633454
rect 547023 633218 571532 633454
rect 571768 633218 571852 633454
rect 572088 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 7876 633134
rect 8112 632898 8196 633134
rect 8432 632898 38032 633134
rect 38268 632898 38352 633134
rect 38588 632898 74032 633134
rect 74268 632898 74352 633134
rect 74588 632898 100443 633134
rect 100679 632898 198919 633134
rect 199155 632898 216399 633134
rect 216635 632898 314875 633134
rect 315111 632898 326032 633134
rect 326268 632898 326352 633134
rect 326588 632898 332355 633134
rect 332591 632898 430831 633134
rect 431067 632898 434032 633134
rect 434268 632898 434352 633134
rect 434588 632898 448311 633134
rect 448547 632898 546787 633134
rect 547023 632898 571532 633134
rect 571768 632898 571852 633134
rect 572088 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 9116 615454
rect 9352 615218 9436 615454
rect 9672 615218 56652 615454
rect 56888 615218 56972 615454
rect 57208 615218 92652 615454
rect 92888 615218 92972 615454
rect 93208 615218 101163 615454
rect 101399 615218 198199 615454
rect 198435 615218 200652 615454
rect 200888 615218 200972 615454
rect 201208 615218 217119 615454
rect 217355 615218 314155 615454
rect 314391 615218 333075 615454
rect 333311 615218 430111 615454
rect 430347 615218 449031 615454
rect 449267 615218 546067 615454
rect 546303 615218 560652 615454
rect 560888 615218 560972 615454
rect 561208 615218 570292 615454
rect 570528 615218 570612 615454
rect 570848 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 9116 615134
rect 9352 614898 9436 615134
rect 9672 614898 56652 615134
rect 56888 614898 56972 615134
rect 57208 614898 92652 615134
rect 92888 614898 92972 615134
rect 93208 614898 101163 615134
rect 101399 614898 198199 615134
rect 198435 614898 200652 615134
rect 200888 614898 200972 615134
rect 201208 614898 217119 615134
rect 217355 614898 314155 615134
rect 314391 614898 333075 615134
rect 333311 614898 430111 615134
rect 430347 614898 449031 615134
rect 449267 614898 546067 615134
rect 546303 614898 560652 615134
rect 560888 614898 560972 615134
rect 561208 614898 570292 615134
rect 570528 614898 570612 615134
rect 570848 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 7876 597454
rect 8112 597218 8196 597454
rect 8432 597218 38032 597454
rect 38268 597218 38352 597454
rect 38588 597218 74032 597454
rect 74268 597218 74352 597454
rect 74588 597218 100443 597454
rect 100679 597218 198919 597454
rect 199155 597218 216399 597454
rect 216635 597218 314875 597454
rect 315111 597218 326032 597454
rect 326268 597218 326352 597454
rect 326588 597218 332355 597454
rect 332591 597218 430831 597454
rect 431067 597218 434032 597454
rect 434268 597218 434352 597454
rect 434588 597218 448311 597454
rect 448547 597218 546787 597454
rect 547023 597218 571532 597454
rect 571768 597218 571852 597454
rect 572088 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 7876 597134
rect 8112 596898 8196 597134
rect 8432 596898 38032 597134
rect 38268 596898 38352 597134
rect 38588 596898 74032 597134
rect 74268 596898 74352 597134
rect 74588 596898 100443 597134
rect 100679 596898 198919 597134
rect 199155 596898 216399 597134
rect 216635 596898 314875 597134
rect 315111 596898 326032 597134
rect 326268 596898 326352 597134
rect 326588 596898 332355 597134
rect 332591 596898 430831 597134
rect 431067 596898 434032 597134
rect 434268 596898 434352 597134
rect 434588 596898 448311 597134
rect 448547 596898 546787 597134
rect 547023 596898 571532 597134
rect 571768 596898 571852 597134
rect 572088 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 9116 579454
rect 9352 579218 9436 579454
rect 9672 579218 56652 579454
rect 56888 579218 56972 579454
rect 57208 579218 92652 579454
rect 92888 579218 92972 579454
rect 93208 579218 128652 579454
rect 128888 579218 128972 579454
rect 129208 579218 164652 579454
rect 164888 579218 164972 579454
rect 165208 579218 200652 579454
rect 200888 579218 200972 579454
rect 201208 579218 236652 579454
rect 236888 579218 236972 579454
rect 237208 579218 272652 579454
rect 272888 579218 272972 579454
rect 273208 579218 308652 579454
rect 308888 579218 308972 579454
rect 309208 579218 344652 579454
rect 344888 579218 344972 579454
rect 345208 579218 380652 579454
rect 380888 579218 380972 579454
rect 381208 579218 416652 579454
rect 416888 579218 416972 579454
rect 417208 579218 452652 579454
rect 452888 579218 452972 579454
rect 453208 579218 488652 579454
rect 488888 579218 488972 579454
rect 489208 579218 524652 579454
rect 524888 579218 524972 579454
rect 525208 579218 560652 579454
rect 560888 579218 560972 579454
rect 561208 579218 570292 579454
rect 570528 579218 570612 579454
rect 570848 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 9116 579134
rect 9352 578898 9436 579134
rect 9672 578898 56652 579134
rect 56888 578898 56972 579134
rect 57208 578898 92652 579134
rect 92888 578898 92972 579134
rect 93208 578898 128652 579134
rect 128888 578898 128972 579134
rect 129208 578898 164652 579134
rect 164888 578898 164972 579134
rect 165208 578898 200652 579134
rect 200888 578898 200972 579134
rect 201208 578898 236652 579134
rect 236888 578898 236972 579134
rect 237208 578898 272652 579134
rect 272888 578898 272972 579134
rect 273208 578898 308652 579134
rect 308888 578898 308972 579134
rect 309208 578898 344652 579134
rect 344888 578898 344972 579134
rect 345208 578898 380652 579134
rect 380888 578898 380972 579134
rect 381208 578898 416652 579134
rect 416888 578898 416972 579134
rect 417208 578898 452652 579134
rect 452888 578898 452972 579134
rect 453208 578898 488652 579134
rect 488888 578898 488972 579134
rect 489208 578898 524652 579134
rect 524888 578898 524972 579134
rect 525208 578898 560652 579134
rect 560888 578898 560972 579134
rect 561208 578898 570292 579134
rect 570528 578898 570612 579134
rect 570848 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 7876 561454
rect 8112 561218 8196 561454
rect 8432 561218 38032 561454
rect 38268 561218 38352 561454
rect 38588 561218 74032 561454
rect 74268 561218 74352 561454
rect 74588 561218 110032 561454
rect 110268 561218 110352 561454
rect 110588 561218 146032 561454
rect 146268 561218 146352 561454
rect 146588 561218 182032 561454
rect 182268 561218 182352 561454
rect 182588 561218 218032 561454
rect 218268 561218 218352 561454
rect 218588 561218 254032 561454
rect 254268 561218 254352 561454
rect 254588 561218 290032 561454
rect 290268 561218 290352 561454
rect 290588 561218 326032 561454
rect 326268 561218 326352 561454
rect 326588 561218 332355 561454
rect 332591 561218 430831 561454
rect 431067 561218 434032 561454
rect 434268 561218 434352 561454
rect 434588 561218 448311 561454
rect 448547 561218 546787 561454
rect 547023 561218 571532 561454
rect 571768 561218 571852 561454
rect 572088 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 7876 561134
rect 8112 560898 8196 561134
rect 8432 560898 38032 561134
rect 38268 560898 38352 561134
rect 38588 560898 74032 561134
rect 74268 560898 74352 561134
rect 74588 560898 110032 561134
rect 110268 560898 110352 561134
rect 110588 560898 146032 561134
rect 146268 560898 146352 561134
rect 146588 560898 182032 561134
rect 182268 560898 182352 561134
rect 182588 560898 218032 561134
rect 218268 560898 218352 561134
rect 218588 560898 254032 561134
rect 254268 560898 254352 561134
rect 254588 560898 290032 561134
rect 290268 560898 290352 561134
rect 290588 560898 326032 561134
rect 326268 560898 326352 561134
rect 326588 560898 332355 561134
rect 332591 560898 430831 561134
rect 431067 560898 434032 561134
rect 434268 560898 434352 561134
rect 434588 560898 448311 561134
rect 448547 560898 546787 561134
rect 547023 560898 571532 561134
rect 571768 560898 571852 561134
rect 572088 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 9116 543454
rect 9352 543218 9436 543454
rect 9672 543218 56652 543454
rect 56888 543218 56972 543454
rect 57208 543218 92652 543454
rect 92888 543218 92972 543454
rect 93208 543218 128652 543454
rect 128888 543218 128972 543454
rect 129208 543218 164652 543454
rect 164888 543218 164972 543454
rect 165208 543218 200652 543454
rect 200888 543218 200972 543454
rect 201208 543218 236652 543454
rect 236888 543218 236972 543454
rect 237208 543218 272652 543454
rect 272888 543218 272972 543454
rect 273208 543218 308652 543454
rect 308888 543218 308972 543454
rect 309208 543218 333075 543454
rect 333311 543218 430111 543454
rect 430347 543218 449031 543454
rect 449267 543218 546067 543454
rect 546303 543218 560652 543454
rect 560888 543218 560972 543454
rect 561208 543218 570292 543454
rect 570528 543218 570612 543454
rect 570848 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 9116 543134
rect 9352 542898 9436 543134
rect 9672 542898 56652 543134
rect 56888 542898 56972 543134
rect 57208 542898 92652 543134
rect 92888 542898 92972 543134
rect 93208 542898 128652 543134
rect 128888 542898 128972 543134
rect 129208 542898 164652 543134
rect 164888 542898 164972 543134
rect 165208 542898 200652 543134
rect 200888 542898 200972 543134
rect 201208 542898 236652 543134
rect 236888 542898 236972 543134
rect 237208 542898 272652 543134
rect 272888 542898 272972 543134
rect 273208 542898 308652 543134
rect 308888 542898 308972 543134
rect 309208 542898 333075 543134
rect 333311 542898 430111 543134
rect 430347 542898 449031 543134
rect 449267 542898 546067 543134
rect 546303 542898 560652 543134
rect 560888 542898 560972 543134
rect 561208 542898 570292 543134
rect 570528 542898 570612 543134
rect 570848 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 7876 525454
rect 8112 525218 8196 525454
rect 8432 525218 38032 525454
rect 38268 525218 38352 525454
rect 38588 525218 74032 525454
rect 74268 525218 74352 525454
rect 74588 525218 110032 525454
rect 110268 525218 110352 525454
rect 110588 525218 146032 525454
rect 146268 525218 146352 525454
rect 146588 525218 182032 525454
rect 182268 525218 182352 525454
rect 182588 525218 218032 525454
rect 218268 525218 218352 525454
rect 218588 525218 254032 525454
rect 254268 525218 254352 525454
rect 254588 525218 290032 525454
rect 290268 525218 290352 525454
rect 290588 525218 326032 525454
rect 326268 525218 326352 525454
rect 326588 525218 332355 525454
rect 332591 525218 430831 525454
rect 431067 525218 434032 525454
rect 434268 525218 434352 525454
rect 434588 525218 448311 525454
rect 448547 525218 546787 525454
rect 547023 525218 571532 525454
rect 571768 525218 571852 525454
rect 572088 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 7876 525134
rect 8112 524898 8196 525134
rect 8432 524898 38032 525134
rect 38268 524898 38352 525134
rect 38588 524898 74032 525134
rect 74268 524898 74352 525134
rect 74588 524898 110032 525134
rect 110268 524898 110352 525134
rect 110588 524898 146032 525134
rect 146268 524898 146352 525134
rect 146588 524898 182032 525134
rect 182268 524898 182352 525134
rect 182588 524898 218032 525134
rect 218268 524898 218352 525134
rect 218588 524898 254032 525134
rect 254268 524898 254352 525134
rect 254588 524898 290032 525134
rect 290268 524898 290352 525134
rect 290588 524898 326032 525134
rect 326268 524898 326352 525134
rect 326588 524898 332355 525134
rect 332591 524898 430831 525134
rect 431067 524898 434032 525134
rect 434268 524898 434352 525134
rect 434588 524898 448311 525134
rect 448547 524898 546787 525134
rect 547023 524898 571532 525134
rect 571768 524898 571852 525134
rect 572088 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 9116 507454
rect 9352 507218 9436 507454
rect 9672 507218 56652 507454
rect 56888 507218 56972 507454
rect 57208 507218 92652 507454
rect 92888 507218 92972 507454
rect 93208 507218 128652 507454
rect 128888 507218 128972 507454
rect 129208 507218 164652 507454
rect 164888 507218 164972 507454
rect 165208 507218 200652 507454
rect 200888 507218 200972 507454
rect 201208 507218 236652 507454
rect 236888 507218 236972 507454
rect 237208 507218 272652 507454
rect 272888 507218 272972 507454
rect 273208 507218 308652 507454
rect 308888 507218 308972 507454
rect 309208 507218 333075 507454
rect 333311 507218 430111 507454
rect 430347 507218 449031 507454
rect 449267 507218 546067 507454
rect 546303 507218 560652 507454
rect 560888 507218 560972 507454
rect 561208 507218 570292 507454
rect 570528 507218 570612 507454
rect 570848 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 9116 507134
rect 9352 506898 9436 507134
rect 9672 506898 56652 507134
rect 56888 506898 56972 507134
rect 57208 506898 92652 507134
rect 92888 506898 92972 507134
rect 93208 506898 128652 507134
rect 128888 506898 128972 507134
rect 129208 506898 164652 507134
rect 164888 506898 164972 507134
rect 165208 506898 200652 507134
rect 200888 506898 200972 507134
rect 201208 506898 236652 507134
rect 236888 506898 236972 507134
rect 237208 506898 272652 507134
rect 272888 506898 272972 507134
rect 273208 506898 308652 507134
rect 308888 506898 308972 507134
rect 309208 506898 333075 507134
rect 333311 506898 430111 507134
rect 430347 506898 449031 507134
rect 449267 506898 546067 507134
rect 546303 506898 560652 507134
rect 560888 506898 560972 507134
rect 561208 506898 570292 507134
rect 570528 506898 570612 507134
rect 570848 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 7876 489454
rect 8112 489218 8196 489454
rect 8432 489218 38032 489454
rect 38268 489218 38352 489454
rect 38588 489218 74032 489454
rect 74268 489218 74352 489454
rect 74588 489218 110032 489454
rect 110268 489218 110352 489454
rect 110588 489218 146032 489454
rect 146268 489218 146352 489454
rect 146588 489218 182032 489454
rect 182268 489218 182352 489454
rect 182588 489218 218032 489454
rect 218268 489218 218352 489454
rect 218588 489218 254032 489454
rect 254268 489218 254352 489454
rect 254588 489218 290032 489454
rect 290268 489218 290352 489454
rect 290588 489218 326032 489454
rect 326268 489218 326352 489454
rect 326588 489218 362032 489454
rect 362268 489218 362352 489454
rect 362588 489218 398032 489454
rect 398268 489218 398352 489454
rect 398588 489218 434032 489454
rect 434268 489218 434352 489454
rect 434588 489218 470032 489454
rect 470268 489218 470352 489454
rect 470588 489218 506032 489454
rect 506268 489218 506352 489454
rect 506588 489218 542032 489454
rect 542268 489218 542352 489454
rect 542588 489218 571532 489454
rect 571768 489218 571852 489454
rect 572088 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 7876 489134
rect 8112 488898 8196 489134
rect 8432 488898 38032 489134
rect 38268 488898 38352 489134
rect 38588 488898 74032 489134
rect 74268 488898 74352 489134
rect 74588 488898 110032 489134
rect 110268 488898 110352 489134
rect 110588 488898 146032 489134
rect 146268 488898 146352 489134
rect 146588 488898 182032 489134
rect 182268 488898 182352 489134
rect 182588 488898 218032 489134
rect 218268 488898 218352 489134
rect 218588 488898 254032 489134
rect 254268 488898 254352 489134
rect 254588 488898 290032 489134
rect 290268 488898 290352 489134
rect 290588 488898 326032 489134
rect 326268 488898 326352 489134
rect 326588 488898 362032 489134
rect 362268 488898 362352 489134
rect 362588 488898 398032 489134
rect 398268 488898 398352 489134
rect 398588 488898 434032 489134
rect 434268 488898 434352 489134
rect 434588 488898 470032 489134
rect 470268 488898 470352 489134
rect 470588 488898 506032 489134
rect 506268 488898 506352 489134
rect 506588 488898 542032 489134
rect 542268 488898 542352 489134
rect 542588 488898 571532 489134
rect 571768 488898 571852 489134
rect 572088 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 9116 471454
rect 9352 471218 9436 471454
rect 9672 471218 56652 471454
rect 56888 471218 56972 471454
rect 57208 471218 92652 471454
rect 92888 471218 92972 471454
rect 93208 471218 128652 471454
rect 128888 471218 128972 471454
rect 129208 471218 164652 471454
rect 164888 471218 164972 471454
rect 165208 471218 200652 471454
rect 200888 471218 200972 471454
rect 201208 471218 236652 471454
rect 236888 471218 236972 471454
rect 237208 471218 272652 471454
rect 272888 471218 272972 471454
rect 273208 471218 308652 471454
rect 308888 471218 308972 471454
rect 309208 471218 333075 471454
rect 333311 471218 430111 471454
rect 430347 471218 449031 471454
rect 449267 471218 546067 471454
rect 546303 471218 560652 471454
rect 560888 471218 560972 471454
rect 561208 471218 570292 471454
rect 570528 471218 570612 471454
rect 570848 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 9116 471134
rect 9352 470898 9436 471134
rect 9672 470898 56652 471134
rect 56888 470898 56972 471134
rect 57208 470898 92652 471134
rect 92888 470898 92972 471134
rect 93208 470898 128652 471134
rect 128888 470898 128972 471134
rect 129208 470898 164652 471134
rect 164888 470898 164972 471134
rect 165208 470898 200652 471134
rect 200888 470898 200972 471134
rect 201208 470898 236652 471134
rect 236888 470898 236972 471134
rect 237208 470898 272652 471134
rect 272888 470898 272972 471134
rect 273208 470898 308652 471134
rect 308888 470898 308972 471134
rect 309208 470898 333075 471134
rect 333311 470898 430111 471134
rect 430347 470898 449031 471134
rect 449267 470898 546067 471134
rect 546303 470898 560652 471134
rect 560888 470898 560972 471134
rect 561208 470898 570292 471134
rect 570528 470898 570612 471134
rect 570848 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 7876 453454
rect 8112 453218 8196 453454
rect 8432 453218 38032 453454
rect 38268 453218 38352 453454
rect 38588 453218 74032 453454
rect 74268 453218 74352 453454
rect 74588 453218 110032 453454
rect 110268 453218 110352 453454
rect 110588 453218 146032 453454
rect 146268 453218 146352 453454
rect 146588 453218 182032 453454
rect 182268 453218 182352 453454
rect 182588 453218 218032 453454
rect 218268 453218 218352 453454
rect 218588 453218 254032 453454
rect 254268 453218 254352 453454
rect 254588 453218 290032 453454
rect 290268 453218 290352 453454
rect 290588 453218 326032 453454
rect 326268 453218 326352 453454
rect 326588 453218 332355 453454
rect 332591 453218 430831 453454
rect 431067 453218 434032 453454
rect 434268 453218 434352 453454
rect 434588 453218 448311 453454
rect 448547 453218 546787 453454
rect 547023 453218 571532 453454
rect 571768 453218 571852 453454
rect 572088 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 7876 453134
rect 8112 452898 8196 453134
rect 8432 452898 38032 453134
rect 38268 452898 38352 453134
rect 38588 452898 74032 453134
rect 74268 452898 74352 453134
rect 74588 452898 110032 453134
rect 110268 452898 110352 453134
rect 110588 452898 146032 453134
rect 146268 452898 146352 453134
rect 146588 452898 182032 453134
rect 182268 452898 182352 453134
rect 182588 452898 218032 453134
rect 218268 452898 218352 453134
rect 218588 452898 254032 453134
rect 254268 452898 254352 453134
rect 254588 452898 290032 453134
rect 290268 452898 290352 453134
rect 290588 452898 326032 453134
rect 326268 452898 326352 453134
rect 326588 452898 332355 453134
rect 332591 452898 430831 453134
rect 431067 452898 434032 453134
rect 434268 452898 434352 453134
rect 434588 452898 448311 453134
rect 448547 452898 546787 453134
rect 547023 452898 571532 453134
rect 571768 452898 571852 453134
rect 572088 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 9116 435454
rect 9352 435218 9436 435454
rect 9672 435218 56652 435454
rect 56888 435218 56972 435454
rect 57208 435218 92652 435454
rect 92888 435218 92972 435454
rect 93208 435218 128652 435454
rect 128888 435218 128972 435454
rect 129208 435218 164652 435454
rect 164888 435218 164972 435454
rect 165208 435218 200652 435454
rect 200888 435218 200972 435454
rect 201208 435218 236652 435454
rect 236888 435218 236972 435454
rect 237208 435218 272652 435454
rect 272888 435218 272972 435454
rect 273208 435218 308652 435454
rect 308888 435218 308972 435454
rect 309208 435218 333075 435454
rect 333311 435218 430111 435454
rect 430347 435218 449031 435454
rect 449267 435218 546067 435454
rect 546303 435218 560652 435454
rect 560888 435218 560972 435454
rect 561208 435218 570292 435454
rect 570528 435218 570612 435454
rect 570848 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 9116 435134
rect 9352 434898 9436 435134
rect 9672 434898 56652 435134
rect 56888 434898 56972 435134
rect 57208 434898 92652 435134
rect 92888 434898 92972 435134
rect 93208 434898 128652 435134
rect 128888 434898 128972 435134
rect 129208 434898 164652 435134
rect 164888 434898 164972 435134
rect 165208 434898 200652 435134
rect 200888 434898 200972 435134
rect 201208 434898 236652 435134
rect 236888 434898 236972 435134
rect 237208 434898 272652 435134
rect 272888 434898 272972 435134
rect 273208 434898 308652 435134
rect 308888 434898 308972 435134
rect 309208 434898 333075 435134
rect 333311 434898 430111 435134
rect 430347 434898 449031 435134
rect 449267 434898 546067 435134
rect 546303 434898 560652 435134
rect 560888 434898 560972 435134
rect 561208 434898 570292 435134
rect 570528 434898 570612 435134
rect 570848 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 7876 417454
rect 8112 417218 8196 417454
rect 8432 417218 38032 417454
rect 38268 417218 38352 417454
rect 38588 417218 74032 417454
rect 74268 417218 74352 417454
rect 74588 417218 110032 417454
rect 110268 417218 110352 417454
rect 110588 417218 146032 417454
rect 146268 417218 146352 417454
rect 146588 417218 182032 417454
rect 182268 417218 182352 417454
rect 182588 417218 218032 417454
rect 218268 417218 218352 417454
rect 218588 417218 254032 417454
rect 254268 417218 254352 417454
rect 254588 417218 290032 417454
rect 290268 417218 290352 417454
rect 290588 417218 326032 417454
rect 326268 417218 326352 417454
rect 326588 417218 332355 417454
rect 332591 417218 430831 417454
rect 431067 417218 434032 417454
rect 434268 417218 434352 417454
rect 434588 417218 448311 417454
rect 448547 417218 546787 417454
rect 547023 417218 571532 417454
rect 571768 417218 571852 417454
rect 572088 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 7876 417134
rect 8112 416898 8196 417134
rect 8432 416898 38032 417134
rect 38268 416898 38352 417134
rect 38588 416898 74032 417134
rect 74268 416898 74352 417134
rect 74588 416898 110032 417134
rect 110268 416898 110352 417134
rect 110588 416898 146032 417134
rect 146268 416898 146352 417134
rect 146588 416898 182032 417134
rect 182268 416898 182352 417134
rect 182588 416898 218032 417134
rect 218268 416898 218352 417134
rect 218588 416898 254032 417134
rect 254268 416898 254352 417134
rect 254588 416898 290032 417134
rect 290268 416898 290352 417134
rect 290588 416898 326032 417134
rect 326268 416898 326352 417134
rect 326588 416898 332355 417134
rect 332591 416898 430831 417134
rect 431067 416898 434032 417134
rect 434268 416898 434352 417134
rect 434588 416898 448311 417134
rect 448547 416898 546787 417134
rect 547023 416898 571532 417134
rect 571768 416898 571852 417134
rect 572088 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 9116 399454
rect 9352 399218 9436 399454
rect 9672 399218 56652 399454
rect 56888 399218 56972 399454
rect 57208 399218 92652 399454
rect 92888 399218 92972 399454
rect 93208 399218 128652 399454
rect 128888 399218 128972 399454
rect 129208 399218 164652 399454
rect 164888 399218 164972 399454
rect 165208 399218 200652 399454
rect 200888 399218 200972 399454
rect 201208 399218 236652 399454
rect 236888 399218 236972 399454
rect 237208 399218 272652 399454
rect 272888 399218 272972 399454
rect 273208 399218 308652 399454
rect 308888 399218 308972 399454
rect 309208 399218 333075 399454
rect 333311 399218 430111 399454
rect 430347 399218 449031 399454
rect 449267 399218 546067 399454
rect 546303 399218 560652 399454
rect 560888 399218 560972 399454
rect 561208 399218 570292 399454
rect 570528 399218 570612 399454
rect 570848 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 9116 399134
rect 9352 398898 9436 399134
rect 9672 398898 56652 399134
rect 56888 398898 56972 399134
rect 57208 398898 92652 399134
rect 92888 398898 92972 399134
rect 93208 398898 128652 399134
rect 128888 398898 128972 399134
rect 129208 398898 164652 399134
rect 164888 398898 164972 399134
rect 165208 398898 200652 399134
rect 200888 398898 200972 399134
rect 201208 398898 236652 399134
rect 236888 398898 236972 399134
rect 237208 398898 272652 399134
rect 272888 398898 272972 399134
rect 273208 398898 308652 399134
rect 308888 398898 308972 399134
rect 309208 398898 333075 399134
rect 333311 398898 430111 399134
rect 430347 398898 449031 399134
rect 449267 398898 546067 399134
rect 546303 398898 560652 399134
rect 560888 398898 560972 399134
rect 561208 398898 570292 399134
rect 570528 398898 570612 399134
rect 570848 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 7876 381454
rect 8112 381218 8196 381454
rect 8432 381218 38032 381454
rect 38268 381218 38352 381454
rect 38588 381218 74032 381454
rect 74268 381218 74352 381454
rect 74588 381218 110032 381454
rect 110268 381218 110352 381454
rect 110588 381218 146032 381454
rect 146268 381218 146352 381454
rect 146588 381218 182032 381454
rect 182268 381218 182352 381454
rect 182588 381218 218032 381454
rect 218268 381218 218352 381454
rect 218588 381218 254032 381454
rect 254268 381218 254352 381454
rect 254588 381218 290032 381454
rect 290268 381218 290352 381454
rect 290588 381218 326032 381454
rect 326268 381218 326352 381454
rect 326588 381218 362032 381454
rect 362268 381218 362352 381454
rect 362588 381218 398032 381454
rect 398268 381218 398352 381454
rect 398588 381218 434032 381454
rect 434268 381218 434352 381454
rect 434588 381218 470032 381454
rect 470268 381218 470352 381454
rect 470588 381218 506032 381454
rect 506268 381218 506352 381454
rect 506588 381218 542032 381454
rect 542268 381218 542352 381454
rect 542588 381218 571532 381454
rect 571768 381218 571852 381454
rect 572088 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 7876 381134
rect 8112 380898 8196 381134
rect 8432 380898 38032 381134
rect 38268 380898 38352 381134
rect 38588 380898 74032 381134
rect 74268 380898 74352 381134
rect 74588 380898 110032 381134
rect 110268 380898 110352 381134
rect 110588 380898 146032 381134
rect 146268 380898 146352 381134
rect 146588 380898 182032 381134
rect 182268 380898 182352 381134
rect 182588 380898 218032 381134
rect 218268 380898 218352 381134
rect 218588 380898 254032 381134
rect 254268 380898 254352 381134
rect 254588 380898 290032 381134
rect 290268 380898 290352 381134
rect 290588 380898 326032 381134
rect 326268 380898 326352 381134
rect 326588 380898 362032 381134
rect 362268 380898 362352 381134
rect 362588 380898 398032 381134
rect 398268 380898 398352 381134
rect 398588 380898 434032 381134
rect 434268 380898 434352 381134
rect 434588 380898 470032 381134
rect 470268 380898 470352 381134
rect 470588 380898 506032 381134
rect 506268 380898 506352 381134
rect 506588 380898 542032 381134
rect 542268 380898 542352 381134
rect 542588 380898 571532 381134
rect 571768 380898 571852 381134
rect 572088 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 9116 363454
rect 9352 363218 9436 363454
rect 9672 363218 56652 363454
rect 56888 363218 56972 363454
rect 57208 363218 92652 363454
rect 92888 363218 92972 363454
rect 93208 363218 128652 363454
rect 128888 363218 128972 363454
rect 129208 363218 164652 363454
rect 164888 363218 164972 363454
rect 165208 363218 200652 363454
rect 200888 363218 200972 363454
rect 201208 363218 236652 363454
rect 236888 363218 236972 363454
rect 237208 363218 272652 363454
rect 272888 363218 272972 363454
rect 273208 363218 308652 363454
rect 308888 363218 308972 363454
rect 309208 363218 333075 363454
rect 333311 363218 430111 363454
rect 430347 363218 449031 363454
rect 449267 363218 546067 363454
rect 546303 363218 560652 363454
rect 560888 363218 560972 363454
rect 561208 363218 570292 363454
rect 570528 363218 570612 363454
rect 570848 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 9116 363134
rect 9352 362898 9436 363134
rect 9672 362898 56652 363134
rect 56888 362898 56972 363134
rect 57208 362898 92652 363134
rect 92888 362898 92972 363134
rect 93208 362898 128652 363134
rect 128888 362898 128972 363134
rect 129208 362898 164652 363134
rect 164888 362898 164972 363134
rect 165208 362898 200652 363134
rect 200888 362898 200972 363134
rect 201208 362898 236652 363134
rect 236888 362898 236972 363134
rect 237208 362898 272652 363134
rect 272888 362898 272972 363134
rect 273208 362898 308652 363134
rect 308888 362898 308972 363134
rect 309208 362898 333075 363134
rect 333311 362898 430111 363134
rect 430347 362898 449031 363134
rect 449267 362898 546067 363134
rect 546303 362898 560652 363134
rect 560888 362898 560972 363134
rect 561208 362898 570292 363134
rect 570528 362898 570612 363134
rect 570848 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 7876 345454
rect 8112 345218 8196 345454
rect 8432 345218 38032 345454
rect 38268 345218 38352 345454
rect 38588 345218 74032 345454
rect 74268 345218 74352 345454
rect 74588 345218 110032 345454
rect 110268 345218 110352 345454
rect 110588 345218 146032 345454
rect 146268 345218 146352 345454
rect 146588 345218 182032 345454
rect 182268 345218 182352 345454
rect 182588 345218 218032 345454
rect 218268 345218 218352 345454
rect 218588 345218 254032 345454
rect 254268 345218 254352 345454
rect 254588 345218 290032 345454
rect 290268 345218 290352 345454
rect 290588 345218 326032 345454
rect 326268 345218 326352 345454
rect 326588 345218 332355 345454
rect 332591 345218 430831 345454
rect 431067 345218 434032 345454
rect 434268 345218 434352 345454
rect 434588 345218 448311 345454
rect 448547 345218 546787 345454
rect 547023 345218 571532 345454
rect 571768 345218 571852 345454
rect 572088 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 7876 345134
rect 8112 344898 8196 345134
rect 8432 344898 38032 345134
rect 38268 344898 38352 345134
rect 38588 344898 74032 345134
rect 74268 344898 74352 345134
rect 74588 344898 110032 345134
rect 110268 344898 110352 345134
rect 110588 344898 146032 345134
rect 146268 344898 146352 345134
rect 146588 344898 182032 345134
rect 182268 344898 182352 345134
rect 182588 344898 218032 345134
rect 218268 344898 218352 345134
rect 218588 344898 254032 345134
rect 254268 344898 254352 345134
rect 254588 344898 290032 345134
rect 290268 344898 290352 345134
rect 290588 344898 326032 345134
rect 326268 344898 326352 345134
rect 326588 344898 332355 345134
rect 332591 344898 430831 345134
rect 431067 344898 434032 345134
rect 434268 344898 434352 345134
rect 434588 344898 448311 345134
rect 448547 344898 546787 345134
rect 547023 344898 571532 345134
rect 571768 344898 571852 345134
rect 572088 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 9116 327454
rect 9352 327218 9436 327454
rect 9672 327218 56652 327454
rect 56888 327218 56972 327454
rect 57208 327218 92652 327454
rect 92888 327218 92972 327454
rect 93208 327218 128652 327454
rect 128888 327218 128972 327454
rect 129208 327218 164652 327454
rect 164888 327218 164972 327454
rect 165208 327218 200652 327454
rect 200888 327218 200972 327454
rect 201208 327218 236652 327454
rect 236888 327218 236972 327454
rect 237208 327218 272652 327454
rect 272888 327218 272972 327454
rect 273208 327218 308652 327454
rect 308888 327218 308972 327454
rect 309208 327218 333075 327454
rect 333311 327218 430111 327454
rect 430347 327218 449031 327454
rect 449267 327218 546067 327454
rect 546303 327218 560652 327454
rect 560888 327218 560972 327454
rect 561208 327218 570292 327454
rect 570528 327218 570612 327454
rect 570848 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 9116 327134
rect 9352 326898 9436 327134
rect 9672 326898 56652 327134
rect 56888 326898 56972 327134
rect 57208 326898 92652 327134
rect 92888 326898 92972 327134
rect 93208 326898 128652 327134
rect 128888 326898 128972 327134
rect 129208 326898 164652 327134
rect 164888 326898 164972 327134
rect 165208 326898 200652 327134
rect 200888 326898 200972 327134
rect 201208 326898 236652 327134
rect 236888 326898 236972 327134
rect 237208 326898 272652 327134
rect 272888 326898 272972 327134
rect 273208 326898 308652 327134
rect 308888 326898 308972 327134
rect 309208 326898 333075 327134
rect 333311 326898 430111 327134
rect 430347 326898 449031 327134
rect 449267 326898 546067 327134
rect 546303 326898 560652 327134
rect 560888 326898 560972 327134
rect 561208 326898 570292 327134
rect 570528 326898 570612 327134
rect 570848 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 7876 309454
rect 8112 309218 8196 309454
rect 8432 309218 38032 309454
rect 38268 309218 38352 309454
rect 38588 309218 74032 309454
rect 74268 309218 74352 309454
rect 74588 309218 110032 309454
rect 110268 309218 110352 309454
rect 110588 309218 146032 309454
rect 146268 309218 146352 309454
rect 146588 309218 182032 309454
rect 182268 309218 182352 309454
rect 182588 309218 218032 309454
rect 218268 309218 218352 309454
rect 218588 309218 254032 309454
rect 254268 309218 254352 309454
rect 254588 309218 290032 309454
rect 290268 309218 290352 309454
rect 290588 309218 326032 309454
rect 326268 309218 326352 309454
rect 326588 309218 332355 309454
rect 332591 309218 430831 309454
rect 431067 309218 434032 309454
rect 434268 309218 434352 309454
rect 434588 309218 448311 309454
rect 448547 309218 546787 309454
rect 547023 309218 571532 309454
rect 571768 309218 571852 309454
rect 572088 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 7876 309134
rect 8112 308898 8196 309134
rect 8432 308898 38032 309134
rect 38268 308898 38352 309134
rect 38588 308898 74032 309134
rect 74268 308898 74352 309134
rect 74588 308898 110032 309134
rect 110268 308898 110352 309134
rect 110588 308898 146032 309134
rect 146268 308898 146352 309134
rect 146588 308898 182032 309134
rect 182268 308898 182352 309134
rect 182588 308898 218032 309134
rect 218268 308898 218352 309134
rect 218588 308898 254032 309134
rect 254268 308898 254352 309134
rect 254588 308898 290032 309134
rect 290268 308898 290352 309134
rect 290588 308898 326032 309134
rect 326268 308898 326352 309134
rect 326588 308898 332355 309134
rect 332591 308898 430831 309134
rect 431067 308898 434032 309134
rect 434268 308898 434352 309134
rect 434588 308898 448311 309134
rect 448547 308898 546787 309134
rect 547023 308898 571532 309134
rect 571768 308898 571852 309134
rect 572088 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 9116 291454
rect 9352 291218 9436 291454
rect 9672 291218 56652 291454
rect 56888 291218 56972 291454
rect 57208 291218 92652 291454
rect 92888 291218 92972 291454
rect 93208 291218 128652 291454
rect 128888 291218 128972 291454
rect 129208 291218 164652 291454
rect 164888 291218 164972 291454
rect 165208 291218 200652 291454
rect 200888 291218 200972 291454
rect 201208 291218 236652 291454
rect 236888 291218 236972 291454
rect 237208 291218 272652 291454
rect 272888 291218 272972 291454
rect 273208 291218 308652 291454
rect 308888 291218 308972 291454
rect 309208 291218 344652 291454
rect 344888 291218 344972 291454
rect 345208 291218 380652 291454
rect 380888 291218 380972 291454
rect 381208 291218 416652 291454
rect 416888 291218 416972 291454
rect 417208 291218 452652 291454
rect 452888 291218 452972 291454
rect 453208 291218 488652 291454
rect 488888 291218 488972 291454
rect 489208 291218 524652 291454
rect 524888 291218 524972 291454
rect 525208 291218 560652 291454
rect 560888 291218 560972 291454
rect 561208 291218 570292 291454
rect 570528 291218 570612 291454
rect 570848 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 9116 291134
rect 9352 290898 9436 291134
rect 9672 290898 56652 291134
rect 56888 290898 56972 291134
rect 57208 290898 92652 291134
rect 92888 290898 92972 291134
rect 93208 290898 128652 291134
rect 128888 290898 128972 291134
rect 129208 290898 164652 291134
rect 164888 290898 164972 291134
rect 165208 290898 200652 291134
rect 200888 290898 200972 291134
rect 201208 290898 236652 291134
rect 236888 290898 236972 291134
rect 237208 290898 272652 291134
rect 272888 290898 272972 291134
rect 273208 290898 308652 291134
rect 308888 290898 308972 291134
rect 309208 290898 344652 291134
rect 344888 290898 344972 291134
rect 345208 290898 380652 291134
rect 380888 290898 380972 291134
rect 381208 290898 416652 291134
rect 416888 290898 416972 291134
rect 417208 290898 452652 291134
rect 452888 290898 452972 291134
rect 453208 290898 488652 291134
rect 488888 290898 488972 291134
rect 489208 290898 524652 291134
rect 524888 290898 524972 291134
rect 525208 290898 560652 291134
rect 560888 290898 560972 291134
rect 561208 290898 570292 291134
rect 570528 290898 570612 291134
rect 570848 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 7876 273454
rect 8112 273218 8196 273454
rect 8432 273218 38032 273454
rect 38268 273218 38352 273454
rect 38588 273218 74032 273454
rect 74268 273218 74352 273454
rect 74588 273218 110032 273454
rect 110268 273218 110352 273454
rect 110588 273218 146032 273454
rect 146268 273218 146352 273454
rect 146588 273218 182032 273454
rect 182268 273218 182352 273454
rect 182588 273218 218032 273454
rect 218268 273218 218352 273454
rect 218588 273218 254032 273454
rect 254268 273218 254352 273454
rect 254588 273218 290032 273454
rect 290268 273218 290352 273454
rect 290588 273218 326032 273454
rect 326268 273218 326352 273454
rect 326588 273218 362032 273454
rect 362268 273218 362352 273454
rect 362588 273218 398032 273454
rect 398268 273218 398352 273454
rect 398588 273218 434032 273454
rect 434268 273218 434352 273454
rect 434588 273218 470032 273454
rect 470268 273218 470352 273454
rect 470588 273218 506032 273454
rect 506268 273218 506352 273454
rect 506588 273218 542032 273454
rect 542268 273218 542352 273454
rect 542588 273218 571532 273454
rect 571768 273218 571852 273454
rect 572088 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 7876 273134
rect 8112 272898 8196 273134
rect 8432 272898 38032 273134
rect 38268 272898 38352 273134
rect 38588 272898 74032 273134
rect 74268 272898 74352 273134
rect 74588 272898 110032 273134
rect 110268 272898 110352 273134
rect 110588 272898 146032 273134
rect 146268 272898 146352 273134
rect 146588 272898 182032 273134
rect 182268 272898 182352 273134
rect 182588 272898 218032 273134
rect 218268 272898 218352 273134
rect 218588 272898 254032 273134
rect 254268 272898 254352 273134
rect 254588 272898 290032 273134
rect 290268 272898 290352 273134
rect 290588 272898 326032 273134
rect 326268 272898 326352 273134
rect 326588 272898 362032 273134
rect 362268 272898 362352 273134
rect 362588 272898 398032 273134
rect 398268 272898 398352 273134
rect 398588 272898 434032 273134
rect 434268 272898 434352 273134
rect 434588 272898 470032 273134
rect 470268 272898 470352 273134
rect 470588 272898 506032 273134
rect 506268 272898 506352 273134
rect 506588 272898 542032 273134
rect 542268 272898 542352 273134
rect 542588 272898 571532 273134
rect 571768 272898 571852 273134
rect 572088 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 9116 255454
rect 9352 255218 9436 255454
rect 9672 255218 56652 255454
rect 56888 255218 56972 255454
rect 57208 255218 92652 255454
rect 92888 255218 92972 255454
rect 93208 255218 128652 255454
rect 128888 255218 128972 255454
rect 129208 255218 164652 255454
rect 164888 255218 164972 255454
rect 165208 255218 200652 255454
rect 200888 255218 200972 255454
rect 201208 255218 236652 255454
rect 236888 255218 236972 255454
rect 237208 255218 272652 255454
rect 272888 255218 272972 255454
rect 273208 255218 308652 255454
rect 308888 255218 308972 255454
rect 309208 255218 344652 255454
rect 344888 255218 344972 255454
rect 345208 255218 380652 255454
rect 380888 255218 380972 255454
rect 381208 255218 416652 255454
rect 416888 255218 416972 255454
rect 417208 255218 452652 255454
rect 452888 255218 452972 255454
rect 453208 255218 488652 255454
rect 488888 255218 488972 255454
rect 489208 255218 524652 255454
rect 524888 255218 524972 255454
rect 525208 255218 560652 255454
rect 560888 255218 560972 255454
rect 561208 255218 570292 255454
rect 570528 255218 570612 255454
rect 570848 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 9116 255134
rect 9352 254898 9436 255134
rect 9672 254898 56652 255134
rect 56888 254898 56972 255134
rect 57208 254898 92652 255134
rect 92888 254898 92972 255134
rect 93208 254898 128652 255134
rect 128888 254898 128972 255134
rect 129208 254898 164652 255134
rect 164888 254898 164972 255134
rect 165208 254898 200652 255134
rect 200888 254898 200972 255134
rect 201208 254898 236652 255134
rect 236888 254898 236972 255134
rect 237208 254898 272652 255134
rect 272888 254898 272972 255134
rect 273208 254898 308652 255134
rect 308888 254898 308972 255134
rect 309208 254898 344652 255134
rect 344888 254898 344972 255134
rect 345208 254898 380652 255134
rect 380888 254898 380972 255134
rect 381208 254898 416652 255134
rect 416888 254898 416972 255134
rect 417208 254898 452652 255134
rect 452888 254898 452972 255134
rect 453208 254898 488652 255134
rect 488888 254898 488972 255134
rect 489208 254898 524652 255134
rect 524888 254898 524972 255134
rect 525208 254898 560652 255134
rect 560888 254898 560972 255134
rect 561208 254898 570292 255134
rect 570528 254898 570612 255134
rect 570848 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 7876 237454
rect 8112 237218 8196 237454
rect 8432 237218 38032 237454
rect 38268 237218 38352 237454
rect 38588 237218 74032 237454
rect 74268 237218 74352 237454
rect 74588 237218 110032 237454
rect 110268 237218 110352 237454
rect 110588 237218 146032 237454
rect 146268 237218 146352 237454
rect 146588 237218 182032 237454
rect 182268 237218 182352 237454
rect 182588 237218 218032 237454
rect 218268 237218 218352 237454
rect 218588 237218 254032 237454
rect 254268 237218 254352 237454
rect 254588 237218 290032 237454
rect 290268 237218 290352 237454
rect 290588 237218 326032 237454
rect 326268 237218 326352 237454
rect 326588 237218 362032 237454
rect 362268 237218 362352 237454
rect 362588 237218 398032 237454
rect 398268 237218 398352 237454
rect 398588 237218 434032 237454
rect 434268 237218 434352 237454
rect 434588 237218 470032 237454
rect 470268 237218 470352 237454
rect 470588 237218 506032 237454
rect 506268 237218 506352 237454
rect 506588 237218 542032 237454
rect 542268 237218 542352 237454
rect 542588 237218 571532 237454
rect 571768 237218 571852 237454
rect 572088 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 7876 237134
rect 8112 236898 8196 237134
rect 8432 236898 38032 237134
rect 38268 236898 38352 237134
rect 38588 236898 74032 237134
rect 74268 236898 74352 237134
rect 74588 236898 110032 237134
rect 110268 236898 110352 237134
rect 110588 236898 146032 237134
rect 146268 236898 146352 237134
rect 146588 236898 182032 237134
rect 182268 236898 182352 237134
rect 182588 236898 218032 237134
rect 218268 236898 218352 237134
rect 218588 236898 254032 237134
rect 254268 236898 254352 237134
rect 254588 236898 290032 237134
rect 290268 236898 290352 237134
rect 290588 236898 326032 237134
rect 326268 236898 326352 237134
rect 326588 236898 362032 237134
rect 362268 236898 362352 237134
rect 362588 236898 398032 237134
rect 398268 236898 398352 237134
rect 398588 236898 434032 237134
rect 434268 236898 434352 237134
rect 434588 236898 470032 237134
rect 470268 236898 470352 237134
rect 470588 236898 506032 237134
rect 506268 236898 506352 237134
rect 506588 236898 542032 237134
rect 542268 236898 542352 237134
rect 542588 236898 571532 237134
rect 571768 236898 571852 237134
rect 572088 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 9116 219454
rect 9352 219218 9436 219454
rect 9672 219218 56652 219454
rect 56888 219218 56972 219454
rect 57208 219218 92652 219454
rect 92888 219218 92972 219454
rect 93208 219218 128652 219454
rect 128888 219218 128972 219454
rect 129208 219218 164652 219454
rect 164888 219218 164972 219454
rect 165208 219218 200652 219454
rect 200888 219218 200972 219454
rect 201208 219218 236652 219454
rect 236888 219218 236972 219454
rect 237208 219218 272652 219454
rect 272888 219218 272972 219454
rect 273208 219218 308652 219454
rect 308888 219218 308972 219454
rect 309208 219218 344652 219454
rect 344888 219218 344972 219454
rect 345208 219218 380652 219454
rect 380888 219218 380972 219454
rect 381208 219218 416652 219454
rect 416888 219218 416972 219454
rect 417208 219218 452652 219454
rect 452888 219218 452972 219454
rect 453208 219218 488652 219454
rect 488888 219218 488972 219454
rect 489208 219218 524652 219454
rect 524888 219218 524972 219454
rect 525208 219218 560652 219454
rect 560888 219218 560972 219454
rect 561208 219218 570292 219454
rect 570528 219218 570612 219454
rect 570848 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 9116 219134
rect 9352 218898 9436 219134
rect 9672 218898 56652 219134
rect 56888 218898 56972 219134
rect 57208 218898 92652 219134
rect 92888 218898 92972 219134
rect 93208 218898 128652 219134
rect 128888 218898 128972 219134
rect 129208 218898 164652 219134
rect 164888 218898 164972 219134
rect 165208 218898 200652 219134
rect 200888 218898 200972 219134
rect 201208 218898 236652 219134
rect 236888 218898 236972 219134
rect 237208 218898 272652 219134
rect 272888 218898 272972 219134
rect 273208 218898 308652 219134
rect 308888 218898 308972 219134
rect 309208 218898 344652 219134
rect 344888 218898 344972 219134
rect 345208 218898 380652 219134
rect 380888 218898 380972 219134
rect 381208 218898 416652 219134
rect 416888 218898 416972 219134
rect 417208 218898 452652 219134
rect 452888 218898 452972 219134
rect 453208 218898 488652 219134
rect 488888 218898 488972 219134
rect 489208 218898 524652 219134
rect 524888 218898 524972 219134
rect 525208 218898 560652 219134
rect 560888 218898 560972 219134
rect 561208 218898 570292 219134
rect 570528 218898 570612 219134
rect 570848 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 7876 201454
rect 8112 201218 8196 201454
rect 8432 201218 38032 201454
rect 38268 201218 38352 201454
rect 38588 201218 74032 201454
rect 74268 201218 74352 201454
rect 74588 201218 110032 201454
rect 110268 201218 110352 201454
rect 110588 201218 146032 201454
rect 146268 201218 146352 201454
rect 146588 201218 182032 201454
rect 182268 201218 182352 201454
rect 182588 201218 218032 201454
rect 218268 201218 218352 201454
rect 218588 201218 254032 201454
rect 254268 201218 254352 201454
rect 254588 201218 290032 201454
rect 290268 201218 290352 201454
rect 290588 201218 326032 201454
rect 326268 201218 326352 201454
rect 326588 201218 362032 201454
rect 362268 201218 362352 201454
rect 362588 201218 398032 201454
rect 398268 201218 398352 201454
rect 398588 201218 434032 201454
rect 434268 201218 434352 201454
rect 434588 201218 470032 201454
rect 470268 201218 470352 201454
rect 470588 201218 506032 201454
rect 506268 201218 506352 201454
rect 506588 201218 542032 201454
rect 542268 201218 542352 201454
rect 542588 201218 571532 201454
rect 571768 201218 571852 201454
rect 572088 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 7876 201134
rect 8112 200898 8196 201134
rect 8432 200898 38032 201134
rect 38268 200898 38352 201134
rect 38588 200898 74032 201134
rect 74268 200898 74352 201134
rect 74588 200898 110032 201134
rect 110268 200898 110352 201134
rect 110588 200898 146032 201134
rect 146268 200898 146352 201134
rect 146588 200898 182032 201134
rect 182268 200898 182352 201134
rect 182588 200898 218032 201134
rect 218268 200898 218352 201134
rect 218588 200898 254032 201134
rect 254268 200898 254352 201134
rect 254588 200898 290032 201134
rect 290268 200898 290352 201134
rect 290588 200898 326032 201134
rect 326268 200898 326352 201134
rect 326588 200898 362032 201134
rect 362268 200898 362352 201134
rect 362588 200898 398032 201134
rect 398268 200898 398352 201134
rect 398588 200898 434032 201134
rect 434268 200898 434352 201134
rect 434588 200898 470032 201134
rect 470268 200898 470352 201134
rect 470588 200898 506032 201134
rect 506268 200898 506352 201134
rect 506588 200898 542032 201134
rect 542268 200898 542352 201134
rect 542588 200898 571532 201134
rect 571768 200898 571852 201134
rect 572088 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 9116 183454
rect 9352 183218 9436 183454
rect 9672 183218 56652 183454
rect 56888 183218 56972 183454
rect 57208 183218 92652 183454
rect 92888 183218 92972 183454
rect 93208 183218 128652 183454
rect 128888 183218 128972 183454
rect 129208 183218 164652 183454
rect 164888 183218 164972 183454
rect 165208 183218 200652 183454
rect 200888 183218 200972 183454
rect 201208 183218 236652 183454
rect 236888 183218 236972 183454
rect 237208 183218 272652 183454
rect 272888 183218 272972 183454
rect 273208 183218 308652 183454
rect 308888 183218 308972 183454
rect 309208 183218 344652 183454
rect 344888 183218 344972 183454
rect 345208 183218 380652 183454
rect 380888 183218 380972 183454
rect 381208 183218 416652 183454
rect 416888 183218 416972 183454
rect 417208 183218 452652 183454
rect 452888 183218 452972 183454
rect 453208 183218 488652 183454
rect 488888 183218 488972 183454
rect 489208 183218 524652 183454
rect 524888 183218 524972 183454
rect 525208 183218 560652 183454
rect 560888 183218 560972 183454
rect 561208 183218 570292 183454
rect 570528 183218 570612 183454
rect 570848 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 9116 183134
rect 9352 182898 9436 183134
rect 9672 182898 56652 183134
rect 56888 182898 56972 183134
rect 57208 182898 92652 183134
rect 92888 182898 92972 183134
rect 93208 182898 128652 183134
rect 128888 182898 128972 183134
rect 129208 182898 164652 183134
rect 164888 182898 164972 183134
rect 165208 182898 200652 183134
rect 200888 182898 200972 183134
rect 201208 182898 236652 183134
rect 236888 182898 236972 183134
rect 237208 182898 272652 183134
rect 272888 182898 272972 183134
rect 273208 182898 308652 183134
rect 308888 182898 308972 183134
rect 309208 182898 344652 183134
rect 344888 182898 344972 183134
rect 345208 182898 380652 183134
rect 380888 182898 380972 183134
rect 381208 182898 416652 183134
rect 416888 182898 416972 183134
rect 417208 182898 452652 183134
rect 452888 182898 452972 183134
rect 453208 182898 488652 183134
rect 488888 182898 488972 183134
rect 489208 182898 524652 183134
rect 524888 182898 524972 183134
rect 525208 182898 560652 183134
rect 560888 182898 560972 183134
rect 561208 182898 570292 183134
rect 570528 182898 570612 183134
rect 570848 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 7876 165454
rect 8112 165218 8196 165454
rect 8432 165218 38032 165454
rect 38268 165218 38352 165454
rect 38588 165218 74032 165454
rect 74268 165218 74352 165454
rect 74588 165218 110032 165454
rect 110268 165218 110352 165454
rect 110588 165218 146032 165454
rect 146268 165218 146352 165454
rect 146588 165218 182032 165454
rect 182268 165218 182352 165454
rect 182588 165218 218032 165454
rect 218268 165218 218352 165454
rect 218588 165218 254032 165454
rect 254268 165218 254352 165454
rect 254588 165218 290032 165454
rect 290268 165218 290352 165454
rect 290588 165218 326032 165454
rect 326268 165218 326352 165454
rect 326588 165218 362032 165454
rect 362268 165218 362352 165454
rect 362588 165218 398032 165454
rect 398268 165218 398352 165454
rect 398588 165218 434032 165454
rect 434268 165218 434352 165454
rect 434588 165218 470032 165454
rect 470268 165218 470352 165454
rect 470588 165218 506032 165454
rect 506268 165218 506352 165454
rect 506588 165218 542032 165454
rect 542268 165218 542352 165454
rect 542588 165218 571532 165454
rect 571768 165218 571852 165454
rect 572088 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 7876 165134
rect 8112 164898 8196 165134
rect 8432 164898 38032 165134
rect 38268 164898 38352 165134
rect 38588 164898 74032 165134
rect 74268 164898 74352 165134
rect 74588 164898 110032 165134
rect 110268 164898 110352 165134
rect 110588 164898 146032 165134
rect 146268 164898 146352 165134
rect 146588 164898 182032 165134
rect 182268 164898 182352 165134
rect 182588 164898 218032 165134
rect 218268 164898 218352 165134
rect 218588 164898 254032 165134
rect 254268 164898 254352 165134
rect 254588 164898 290032 165134
rect 290268 164898 290352 165134
rect 290588 164898 326032 165134
rect 326268 164898 326352 165134
rect 326588 164898 362032 165134
rect 362268 164898 362352 165134
rect 362588 164898 398032 165134
rect 398268 164898 398352 165134
rect 398588 164898 434032 165134
rect 434268 164898 434352 165134
rect 434588 164898 470032 165134
rect 470268 164898 470352 165134
rect 470588 164898 506032 165134
rect 506268 164898 506352 165134
rect 506588 164898 542032 165134
rect 542268 164898 542352 165134
rect 542588 164898 571532 165134
rect 571768 164898 571852 165134
rect 572088 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 9116 147454
rect 9352 147218 9436 147454
rect 9672 147218 56652 147454
rect 56888 147218 56972 147454
rect 57208 147218 92652 147454
rect 92888 147218 92972 147454
rect 93208 147218 128652 147454
rect 128888 147218 128972 147454
rect 129208 147218 164652 147454
rect 164888 147218 164972 147454
rect 165208 147218 200652 147454
rect 200888 147218 200972 147454
rect 201208 147218 236652 147454
rect 236888 147218 236972 147454
rect 237208 147218 272652 147454
rect 272888 147218 272972 147454
rect 273208 147218 308652 147454
rect 308888 147218 308972 147454
rect 309208 147218 344652 147454
rect 344888 147218 344972 147454
rect 345208 147218 380652 147454
rect 380888 147218 380972 147454
rect 381208 147218 416652 147454
rect 416888 147218 416972 147454
rect 417208 147218 452652 147454
rect 452888 147218 452972 147454
rect 453208 147218 488652 147454
rect 488888 147218 488972 147454
rect 489208 147218 524652 147454
rect 524888 147218 524972 147454
rect 525208 147218 560652 147454
rect 560888 147218 560972 147454
rect 561208 147218 570292 147454
rect 570528 147218 570612 147454
rect 570848 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 9116 147134
rect 9352 146898 9436 147134
rect 9672 146898 56652 147134
rect 56888 146898 56972 147134
rect 57208 146898 92652 147134
rect 92888 146898 92972 147134
rect 93208 146898 128652 147134
rect 128888 146898 128972 147134
rect 129208 146898 164652 147134
rect 164888 146898 164972 147134
rect 165208 146898 200652 147134
rect 200888 146898 200972 147134
rect 201208 146898 236652 147134
rect 236888 146898 236972 147134
rect 237208 146898 272652 147134
rect 272888 146898 272972 147134
rect 273208 146898 308652 147134
rect 308888 146898 308972 147134
rect 309208 146898 344652 147134
rect 344888 146898 344972 147134
rect 345208 146898 380652 147134
rect 380888 146898 380972 147134
rect 381208 146898 416652 147134
rect 416888 146898 416972 147134
rect 417208 146898 452652 147134
rect 452888 146898 452972 147134
rect 453208 146898 488652 147134
rect 488888 146898 488972 147134
rect 489208 146898 524652 147134
rect 524888 146898 524972 147134
rect 525208 146898 560652 147134
rect 560888 146898 560972 147134
rect 561208 146898 570292 147134
rect 570528 146898 570612 147134
rect 570848 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 7876 129454
rect 8112 129218 8196 129454
rect 8432 129218 38032 129454
rect 38268 129218 38352 129454
rect 38588 129218 74032 129454
rect 74268 129218 74352 129454
rect 74588 129218 110032 129454
rect 110268 129218 110352 129454
rect 110588 129218 146032 129454
rect 146268 129218 146352 129454
rect 146588 129218 182032 129454
rect 182268 129218 182352 129454
rect 182588 129218 218032 129454
rect 218268 129218 218352 129454
rect 218588 129218 254032 129454
rect 254268 129218 254352 129454
rect 254588 129218 290032 129454
rect 290268 129218 290352 129454
rect 290588 129218 326032 129454
rect 326268 129218 326352 129454
rect 326588 129218 362032 129454
rect 362268 129218 362352 129454
rect 362588 129218 398032 129454
rect 398268 129218 398352 129454
rect 398588 129218 434032 129454
rect 434268 129218 434352 129454
rect 434588 129218 470032 129454
rect 470268 129218 470352 129454
rect 470588 129218 506032 129454
rect 506268 129218 506352 129454
rect 506588 129218 542032 129454
rect 542268 129218 542352 129454
rect 542588 129218 571532 129454
rect 571768 129218 571852 129454
rect 572088 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 7876 129134
rect 8112 128898 8196 129134
rect 8432 128898 38032 129134
rect 38268 128898 38352 129134
rect 38588 128898 74032 129134
rect 74268 128898 74352 129134
rect 74588 128898 110032 129134
rect 110268 128898 110352 129134
rect 110588 128898 146032 129134
rect 146268 128898 146352 129134
rect 146588 128898 182032 129134
rect 182268 128898 182352 129134
rect 182588 128898 218032 129134
rect 218268 128898 218352 129134
rect 218588 128898 254032 129134
rect 254268 128898 254352 129134
rect 254588 128898 290032 129134
rect 290268 128898 290352 129134
rect 290588 128898 326032 129134
rect 326268 128898 326352 129134
rect 326588 128898 362032 129134
rect 362268 128898 362352 129134
rect 362588 128898 398032 129134
rect 398268 128898 398352 129134
rect 398588 128898 434032 129134
rect 434268 128898 434352 129134
rect 434588 128898 470032 129134
rect 470268 128898 470352 129134
rect 470588 128898 506032 129134
rect 506268 128898 506352 129134
rect 506588 128898 542032 129134
rect 542268 128898 542352 129134
rect 542588 128898 571532 129134
rect 571768 128898 571852 129134
rect 572088 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 9116 111454
rect 9352 111218 9436 111454
rect 9672 111218 56652 111454
rect 56888 111218 56972 111454
rect 57208 111218 92652 111454
rect 92888 111218 92972 111454
rect 93208 111218 128652 111454
rect 128888 111218 128972 111454
rect 129208 111218 164652 111454
rect 164888 111218 164972 111454
rect 165208 111218 200652 111454
rect 200888 111218 200972 111454
rect 201208 111218 236652 111454
rect 236888 111218 236972 111454
rect 237208 111218 272652 111454
rect 272888 111218 272972 111454
rect 273208 111218 308652 111454
rect 308888 111218 308972 111454
rect 309208 111218 344652 111454
rect 344888 111218 344972 111454
rect 345208 111218 380652 111454
rect 380888 111218 380972 111454
rect 381208 111218 416652 111454
rect 416888 111218 416972 111454
rect 417208 111218 452652 111454
rect 452888 111218 452972 111454
rect 453208 111218 488652 111454
rect 488888 111218 488972 111454
rect 489208 111218 524652 111454
rect 524888 111218 524972 111454
rect 525208 111218 560652 111454
rect 560888 111218 560972 111454
rect 561208 111218 570292 111454
rect 570528 111218 570612 111454
rect 570848 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 9116 111134
rect 9352 110898 9436 111134
rect 9672 110898 56652 111134
rect 56888 110898 56972 111134
rect 57208 110898 92652 111134
rect 92888 110898 92972 111134
rect 93208 110898 128652 111134
rect 128888 110898 128972 111134
rect 129208 110898 164652 111134
rect 164888 110898 164972 111134
rect 165208 110898 200652 111134
rect 200888 110898 200972 111134
rect 201208 110898 236652 111134
rect 236888 110898 236972 111134
rect 237208 110898 272652 111134
rect 272888 110898 272972 111134
rect 273208 110898 308652 111134
rect 308888 110898 308972 111134
rect 309208 110898 344652 111134
rect 344888 110898 344972 111134
rect 345208 110898 380652 111134
rect 380888 110898 380972 111134
rect 381208 110898 416652 111134
rect 416888 110898 416972 111134
rect 417208 110898 452652 111134
rect 452888 110898 452972 111134
rect 453208 110898 488652 111134
rect 488888 110898 488972 111134
rect 489208 110898 524652 111134
rect 524888 110898 524972 111134
rect 525208 110898 560652 111134
rect 560888 110898 560972 111134
rect 561208 110898 570292 111134
rect 570528 110898 570612 111134
rect 570848 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 7876 93454
rect 8112 93218 8196 93454
rect 8432 93218 38032 93454
rect 38268 93218 38352 93454
rect 38588 93218 74032 93454
rect 74268 93218 74352 93454
rect 74588 93218 110032 93454
rect 110268 93218 110352 93454
rect 110588 93218 146032 93454
rect 146268 93218 146352 93454
rect 146588 93218 182032 93454
rect 182268 93218 182352 93454
rect 182588 93218 218032 93454
rect 218268 93218 218352 93454
rect 218588 93218 254032 93454
rect 254268 93218 254352 93454
rect 254588 93218 290032 93454
rect 290268 93218 290352 93454
rect 290588 93218 326032 93454
rect 326268 93218 326352 93454
rect 326588 93218 362032 93454
rect 362268 93218 362352 93454
rect 362588 93218 398032 93454
rect 398268 93218 398352 93454
rect 398588 93218 434032 93454
rect 434268 93218 434352 93454
rect 434588 93218 470032 93454
rect 470268 93218 470352 93454
rect 470588 93218 506032 93454
rect 506268 93218 506352 93454
rect 506588 93218 542032 93454
rect 542268 93218 542352 93454
rect 542588 93218 571532 93454
rect 571768 93218 571852 93454
rect 572088 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 7876 93134
rect 8112 92898 8196 93134
rect 8432 92898 38032 93134
rect 38268 92898 38352 93134
rect 38588 92898 74032 93134
rect 74268 92898 74352 93134
rect 74588 92898 110032 93134
rect 110268 92898 110352 93134
rect 110588 92898 146032 93134
rect 146268 92898 146352 93134
rect 146588 92898 182032 93134
rect 182268 92898 182352 93134
rect 182588 92898 218032 93134
rect 218268 92898 218352 93134
rect 218588 92898 254032 93134
rect 254268 92898 254352 93134
rect 254588 92898 290032 93134
rect 290268 92898 290352 93134
rect 290588 92898 326032 93134
rect 326268 92898 326352 93134
rect 326588 92898 362032 93134
rect 362268 92898 362352 93134
rect 362588 92898 398032 93134
rect 398268 92898 398352 93134
rect 398588 92898 434032 93134
rect 434268 92898 434352 93134
rect 434588 92898 470032 93134
rect 470268 92898 470352 93134
rect 470588 92898 506032 93134
rect 506268 92898 506352 93134
rect 506588 92898 542032 93134
rect 542268 92898 542352 93134
rect 542588 92898 571532 93134
rect 571768 92898 571852 93134
rect 572088 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 9116 75454
rect 9352 75218 9436 75454
rect 9672 75218 56652 75454
rect 56888 75218 56972 75454
rect 57208 75218 92652 75454
rect 92888 75218 92972 75454
rect 93208 75218 128652 75454
rect 128888 75218 128972 75454
rect 129208 75218 164652 75454
rect 164888 75218 164972 75454
rect 165208 75218 200652 75454
rect 200888 75218 200972 75454
rect 201208 75218 236652 75454
rect 236888 75218 236972 75454
rect 237208 75218 272652 75454
rect 272888 75218 272972 75454
rect 273208 75218 308652 75454
rect 308888 75218 308972 75454
rect 309208 75218 344652 75454
rect 344888 75218 344972 75454
rect 345208 75218 380652 75454
rect 380888 75218 380972 75454
rect 381208 75218 416652 75454
rect 416888 75218 416972 75454
rect 417208 75218 452652 75454
rect 452888 75218 452972 75454
rect 453208 75218 488652 75454
rect 488888 75218 488972 75454
rect 489208 75218 524652 75454
rect 524888 75218 524972 75454
rect 525208 75218 560652 75454
rect 560888 75218 560972 75454
rect 561208 75218 570292 75454
rect 570528 75218 570612 75454
rect 570848 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 9116 75134
rect 9352 74898 9436 75134
rect 9672 74898 56652 75134
rect 56888 74898 56972 75134
rect 57208 74898 92652 75134
rect 92888 74898 92972 75134
rect 93208 74898 128652 75134
rect 128888 74898 128972 75134
rect 129208 74898 164652 75134
rect 164888 74898 164972 75134
rect 165208 74898 200652 75134
rect 200888 74898 200972 75134
rect 201208 74898 236652 75134
rect 236888 74898 236972 75134
rect 237208 74898 272652 75134
rect 272888 74898 272972 75134
rect 273208 74898 308652 75134
rect 308888 74898 308972 75134
rect 309208 74898 344652 75134
rect 344888 74898 344972 75134
rect 345208 74898 380652 75134
rect 380888 74898 380972 75134
rect 381208 74898 416652 75134
rect 416888 74898 416972 75134
rect 417208 74898 452652 75134
rect 452888 74898 452972 75134
rect 453208 74898 488652 75134
rect 488888 74898 488972 75134
rect 489208 74898 524652 75134
rect 524888 74898 524972 75134
rect 525208 74898 560652 75134
rect 560888 74898 560972 75134
rect 561208 74898 570292 75134
rect 570528 74898 570612 75134
rect 570848 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 7876 57454
rect 8112 57218 8196 57454
rect 8432 57218 38032 57454
rect 38268 57218 38352 57454
rect 38588 57218 74032 57454
rect 74268 57218 74352 57454
rect 74588 57218 110032 57454
rect 110268 57218 110352 57454
rect 110588 57218 146032 57454
rect 146268 57218 146352 57454
rect 146588 57218 182032 57454
rect 182268 57218 182352 57454
rect 182588 57218 218032 57454
rect 218268 57218 218352 57454
rect 218588 57218 254032 57454
rect 254268 57218 254352 57454
rect 254588 57218 290032 57454
rect 290268 57218 290352 57454
rect 290588 57218 326032 57454
rect 326268 57218 326352 57454
rect 326588 57218 362032 57454
rect 362268 57218 362352 57454
rect 362588 57218 398032 57454
rect 398268 57218 398352 57454
rect 398588 57218 434032 57454
rect 434268 57218 434352 57454
rect 434588 57218 470032 57454
rect 470268 57218 470352 57454
rect 470588 57218 506032 57454
rect 506268 57218 506352 57454
rect 506588 57218 542032 57454
rect 542268 57218 542352 57454
rect 542588 57218 571532 57454
rect 571768 57218 571852 57454
rect 572088 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 7876 57134
rect 8112 56898 8196 57134
rect 8432 56898 38032 57134
rect 38268 56898 38352 57134
rect 38588 56898 74032 57134
rect 74268 56898 74352 57134
rect 74588 56898 110032 57134
rect 110268 56898 110352 57134
rect 110588 56898 146032 57134
rect 146268 56898 146352 57134
rect 146588 56898 182032 57134
rect 182268 56898 182352 57134
rect 182588 56898 218032 57134
rect 218268 56898 218352 57134
rect 218588 56898 254032 57134
rect 254268 56898 254352 57134
rect 254588 56898 290032 57134
rect 290268 56898 290352 57134
rect 290588 56898 326032 57134
rect 326268 56898 326352 57134
rect 326588 56898 362032 57134
rect 362268 56898 362352 57134
rect 362588 56898 398032 57134
rect 398268 56898 398352 57134
rect 398588 56898 434032 57134
rect 434268 56898 434352 57134
rect 434588 56898 470032 57134
rect 470268 56898 470352 57134
rect 470588 56898 506032 57134
rect 506268 56898 506352 57134
rect 506588 56898 542032 57134
rect 542268 56898 542352 57134
rect 542588 56898 571532 57134
rect 571768 56898 571852 57134
rect 572088 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 9116 39454
rect 9352 39218 9436 39454
rect 9672 39218 56652 39454
rect 56888 39218 56972 39454
rect 57208 39218 92652 39454
rect 92888 39218 92972 39454
rect 93208 39218 128652 39454
rect 128888 39218 128972 39454
rect 129208 39218 164652 39454
rect 164888 39218 164972 39454
rect 165208 39218 200652 39454
rect 200888 39218 200972 39454
rect 201208 39218 236652 39454
rect 236888 39218 236972 39454
rect 237208 39218 272652 39454
rect 272888 39218 272972 39454
rect 273208 39218 308652 39454
rect 308888 39218 308972 39454
rect 309208 39218 344652 39454
rect 344888 39218 344972 39454
rect 345208 39218 380652 39454
rect 380888 39218 380972 39454
rect 381208 39218 416652 39454
rect 416888 39218 416972 39454
rect 417208 39218 452652 39454
rect 452888 39218 452972 39454
rect 453208 39218 488652 39454
rect 488888 39218 488972 39454
rect 489208 39218 524652 39454
rect 524888 39218 524972 39454
rect 525208 39218 560652 39454
rect 560888 39218 560972 39454
rect 561208 39218 570292 39454
rect 570528 39218 570612 39454
rect 570848 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 9116 39134
rect 9352 38898 9436 39134
rect 9672 38898 56652 39134
rect 56888 38898 56972 39134
rect 57208 38898 92652 39134
rect 92888 38898 92972 39134
rect 93208 38898 128652 39134
rect 128888 38898 128972 39134
rect 129208 38898 164652 39134
rect 164888 38898 164972 39134
rect 165208 38898 200652 39134
rect 200888 38898 200972 39134
rect 201208 38898 236652 39134
rect 236888 38898 236972 39134
rect 237208 38898 272652 39134
rect 272888 38898 272972 39134
rect 273208 38898 308652 39134
rect 308888 38898 308972 39134
rect 309208 38898 344652 39134
rect 344888 38898 344972 39134
rect 345208 38898 380652 39134
rect 380888 38898 380972 39134
rect 381208 38898 416652 39134
rect 416888 38898 416972 39134
rect 417208 38898 452652 39134
rect 452888 38898 452972 39134
rect 453208 38898 488652 39134
rect 488888 38898 488972 39134
rect 489208 38898 524652 39134
rect 524888 38898 524972 39134
rect 525208 38898 560652 39134
rect 560888 38898 560972 39134
rect 561208 38898 570292 39134
rect 570528 38898 570612 39134
rect 570848 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 7876 21454
rect 8112 21218 8196 21454
rect 8432 21218 38032 21454
rect 38268 21218 38352 21454
rect 38588 21218 74032 21454
rect 74268 21218 74352 21454
rect 74588 21218 110032 21454
rect 110268 21218 110352 21454
rect 110588 21218 146032 21454
rect 146268 21218 146352 21454
rect 146588 21218 182032 21454
rect 182268 21218 182352 21454
rect 182588 21218 218032 21454
rect 218268 21218 218352 21454
rect 218588 21218 254032 21454
rect 254268 21218 254352 21454
rect 254588 21218 290032 21454
rect 290268 21218 290352 21454
rect 290588 21218 326032 21454
rect 326268 21218 326352 21454
rect 326588 21218 362032 21454
rect 362268 21218 362352 21454
rect 362588 21218 398032 21454
rect 398268 21218 398352 21454
rect 398588 21218 434032 21454
rect 434268 21218 434352 21454
rect 434588 21218 470032 21454
rect 470268 21218 470352 21454
rect 470588 21218 506032 21454
rect 506268 21218 506352 21454
rect 506588 21218 542032 21454
rect 542268 21218 542352 21454
rect 542588 21218 571532 21454
rect 571768 21218 571852 21454
rect 572088 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 7876 21134
rect 8112 20898 8196 21134
rect 8432 20898 38032 21134
rect 38268 20898 38352 21134
rect 38588 20898 74032 21134
rect 74268 20898 74352 21134
rect 74588 20898 110032 21134
rect 110268 20898 110352 21134
rect 110588 20898 146032 21134
rect 146268 20898 146352 21134
rect 146588 20898 182032 21134
rect 182268 20898 182352 21134
rect 182588 20898 218032 21134
rect 218268 20898 218352 21134
rect 218588 20898 254032 21134
rect 254268 20898 254352 21134
rect 254588 20898 290032 21134
rect 290268 20898 290352 21134
rect 290588 20898 326032 21134
rect 326268 20898 326352 21134
rect 326588 20898 362032 21134
rect 362268 20898 362352 21134
rect 362588 20898 398032 21134
rect 398268 20898 398352 21134
rect 398588 20898 434032 21134
rect 434268 20898 434352 21134
rect 434588 20898 470032 21134
rect 470268 20898 470352 21134
rect 470588 20898 506032 21134
rect 506268 20898 506352 21134
rect 506588 20898 542032 21134
rect 542268 20898 542352 21134
rect 542588 20898 571532 21134
rect 571768 20898 571852 21134
rect 572088 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 0
transform 1 0 4000 0 1 4000
box 0 0 571964 694008
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 700008 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 700008 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 700008 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 700008 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 700008 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 700008 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 700008 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 700008 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 700008 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 700008 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 700008 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 700008 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 700008 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 700008 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 700008 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 700008 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 700008 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 700008 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 700008 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 700008 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 700008 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 700008 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 700008 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 700008 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 700008 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 700008 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 700008 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 700008 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 700008 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 700008 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 700008 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 700008 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 700008 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 700008 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 700008 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 700008 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 700008 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 700008 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 700008 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 700008 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 700008 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 700008 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 700008 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 700008 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 700008 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 700008 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 700008 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 700008 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 700008 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 700008 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 700008 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 700008 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 700008 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 700008 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 700008 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 700008 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 700008 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 700008 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 700008 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 700008 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 700008 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 700008 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 700008 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 700008 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 700008 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 700008 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 700008 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 700008 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 700008 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 700008 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 700008 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 700008 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 700008 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 700008 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 700008 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 700008 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 700008 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 700008 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 700008 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 700008 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 700008 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 700008 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 700008 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 700008 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 700008 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 700008 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 700008 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 700008 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 700008 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 700008 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 700008 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 700008 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 700008 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 700008 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 700008 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 700008 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 700008 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 700008 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 700008 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 700008 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 700008 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 700008 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 700008 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 700008 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 700008 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 700008 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 700008 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 700008 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 700008 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 700008 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 700008 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 700008 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 700008 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 700008 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 700008 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 700008 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 700008 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 700008 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 700008 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 700008 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 700008 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 700008 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 700008 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 700008 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 700008 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 700008 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 700008 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 700008 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 700008 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
