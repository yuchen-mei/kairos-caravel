magic
tech sky130A
timestamp 1656789359
<< obsli1 >>
rect 2000 2000 287982 349004
<< obsm1 >>
rect 283 4 291817 350400
<< metal2 >>
rect 4043 351760 4099 352480
rect 12139 351760 12195 352480
rect 20235 351760 20291 352480
rect 28377 351760 28433 352480
rect 36473 351760 36529 352480
rect 44569 351760 44625 352480
rect 52711 351760 52767 352480
rect 60807 351760 60863 352480
rect 68903 351760 68959 352480
rect 77045 351760 77101 352480
rect 85141 351760 85197 352480
rect 93237 351760 93293 352480
rect 101379 351760 101435 352480
rect 109475 351760 109531 352480
rect 117571 351760 117627 352480
rect 125713 351760 125769 352480
rect 133809 351760 133865 352480
rect 141905 351760 141961 352480
rect 150047 351760 150103 352480
rect 158143 351760 158199 352480
rect 166239 351760 166295 352480
rect 174381 351760 174437 352480
rect 182477 351760 182533 352480
rect 190573 351760 190629 352480
rect 198715 351760 198771 352480
rect 206811 351760 206867 352480
rect 214907 351760 214963 352480
rect 223049 351760 223105 352480
rect 231145 351760 231201 352480
rect 239241 351760 239297 352480
rect 247383 351760 247439 352480
rect 255479 351760 255535 352480
rect 263575 351760 263631 352480
rect 271717 351760 271773 352480
rect 279813 351760 279869 352480
rect 287909 351760 287965 352480
rect 271 -480 327 240
rect 823 -480 879 240
rect 1421 -480 1477 240
rect 2019 -480 2075 240
rect 2617 -480 2673 240
rect 3215 -480 3271 240
rect 3813 -480 3869 240
rect 4365 -480 4421 240
rect 4963 -480 5019 240
rect 5561 -480 5617 240
rect 6159 -480 6215 240
rect 6757 -480 6813 240
rect 7355 -480 7411 240
rect 7953 -480 8009 240
rect 8505 -480 8561 240
rect 9103 -480 9159 240
rect 9701 -480 9757 240
rect 10299 -480 10355 240
rect 10897 -480 10953 240
rect 11495 -480 11551 240
rect 12093 -480 12149 240
rect 12645 -480 12701 240
rect 13243 -480 13299 240
rect 13841 -480 13897 240
rect 14439 -480 14495 240
rect 15037 -480 15093 240
rect 15635 -480 15691 240
rect 16187 -480 16243 240
rect 16785 -480 16841 240
rect 17383 -480 17439 240
rect 17981 -480 18037 240
rect 18579 -480 18635 240
rect 19177 -480 19233 240
rect 19775 -480 19831 240
rect 20327 -480 20383 240
rect 20925 -480 20981 240
rect 21523 -480 21579 240
rect 22121 -480 22177 240
rect 22719 -480 22775 240
rect 23317 -480 23373 240
rect 23915 -480 23971 240
rect 24467 -480 24523 240
rect 25065 -480 25121 240
rect 25663 -480 25719 240
rect 26261 -480 26317 240
rect 26859 -480 26915 240
rect 27457 -480 27513 240
rect 28009 -480 28065 240
rect 28607 -480 28663 240
rect 29205 -480 29261 240
rect 29803 -480 29859 240
rect 30401 -480 30457 240
rect 30999 -480 31055 240
rect 31597 -480 31653 240
rect 32149 -480 32205 240
rect 32747 -480 32803 240
rect 33345 -480 33401 240
rect 33943 -480 33999 240
rect 34541 -480 34597 240
rect 35139 -480 35195 240
rect 35737 -480 35793 240
rect 36289 -480 36345 240
rect 36887 -480 36943 240
rect 37485 -480 37541 240
rect 38083 -480 38139 240
rect 38681 -480 38737 240
rect 39279 -480 39335 240
rect 39831 -480 39887 240
rect 40429 -480 40485 240
rect 41027 -480 41083 240
rect 41625 -480 41681 240
rect 42223 -480 42279 240
rect 42821 -480 42877 240
rect 43419 -480 43475 240
rect 43971 -480 44027 240
rect 44569 -480 44625 240
rect 45167 -480 45223 240
rect 45765 -480 45821 240
rect 46363 -480 46419 240
rect 46961 -480 47017 240
rect 47559 -480 47615 240
rect 48111 -480 48167 240
rect 48709 -480 48765 240
rect 49307 -480 49363 240
rect 49905 -480 49961 240
rect 50503 -480 50559 240
rect 51101 -480 51157 240
rect 51653 -480 51709 240
rect 52251 -480 52307 240
rect 52849 -480 52905 240
rect 53447 -480 53503 240
rect 54045 -480 54101 240
rect 54643 -480 54699 240
rect 55241 -480 55297 240
rect 55793 -480 55849 240
rect 56391 -480 56447 240
rect 56989 -480 57045 240
rect 57587 -480 57643 240
rect 58185 -480 58241 240
rect 58783 -480 58839 240
rect 59381 -480 59437 240
rect 59933 -480 59989 240
rect 60531 -480 60587 240
rect 61129 -480 61185 240
rect 61727 -480 61783 240
rect 62325 -480 62381 240
rect 62923 -480 62979 240
rect 63475 -480 63531 240
rect 64073 -480 64129 240
rect 64671 -480 64727 240
rect 65269 -480 65325 240
rect 65867 -480 65923 240
rect 66465 -480 66521 240
rect 67063 -480 67119 240
rect 67615 -480 67671 240
rect 68213 -480 68269 240
rect 68811 -480 68867 240
rect 69409 -480 69465 240
rect 70007 -480 70063 240
rect 70605 -480 70661 240
rect 71203 -480 71259 240
rect 71755 -480 71811 240
rect 72353 -480 72409 240
rect 72951 -480 73007 240
rect 73549 -480 73605 240
rect 74147 -480 74203 240
rect 74745 -480 74801 240
rect 75297 -480 75353 240
rect 75895 -480 75951 240
rect 76493 -480 76549 240
rect 77091 -480 77147 240
rect 77689 -480 77745 240
rect 78287 -480 78343 240
rect 78885 -480 78941 240
rect 79437 -480 79493 240
rect 80035 -480 80091 240
rect 80633 -480 80689 240
rect 81231 -480 81287 240
rect 81829 -480 81885 240
rect 82427 -480 82483 240
rect 83025 -480 83081 240
rect 83577 -480 83633 240
rect 84175 -480 84231 240
rect 84773 -480 84829 240
rect 85371 -480 85427 240
rect 85969 -480 86025 240
rect 86567 -480 86623 240
rect 87119 -480 87175 240
rect 87717 -480 87773 240
rect 88315 -480 88371 240
rect 88913 -480 88969 240
rect 89511 -480 89567 240
rect 90109 -480 90165 240
rect 90707 -480 90763 240
rect 91259 -480 91315 240
rect 91857 -480 91913 240
rect 92455 -480 92511 240
rect 93053 -480 93109 240
rect 93651 -480 93707 240
rect 94249 -480 94305 240
rect 94847 -480 94903 240
rect 95399 -480 95455 240
rect 95997 -480 96053 240
rect 96595 -480 96651 240
rect 97193 -480 97249 240
rect 97791 -480 97847 240
rect 98389 -480 98445 240
rect 98941 -480 98997 240
rect 99539 -480 99595 240
rect 100137 -480 100193 240
rect 100735 -480 100791 240
rect 101333 -480 101389 240
rect 101931 -480 101987 240
rect 102529 -480 102585 240
rect 103081 -480 103137 240
rect 103679 -480 103735 240
rect 104277 -480 104333 240
rect 104875 -480 104931 240
rect 105473 -480 105529 240
rect 106071 -480 106127 240
rect 106669 -480 106725 240
rect 107221 -480 107277 240
rect 107819 -480 107875 240
rect 108417 -480 108473 240
rect 109015 -480 109071 240
rect 109613 -480 109669 240
rect 110211 -480 110267 240
rect 110763 -480 110819 240
rect 111361 -480 111417 240
rect 111959 -480 112015 240
rect 112557 -480 112613 240
rect 113155 -480 113211 240
rect 113753 -480 113809 240
rect 114351 -480 114407 240
rect 114903 -480 114959 240
rect 115501 -480 115557 240
rect 116099 -480 116155 240
rect 116697 -480 116753 240
rect 117295 -480 117351 240
rect 117893 -480 117949 240
rect 118491 -480 118547 240
rect 119043 -480 119099 240
rect 119641 -480 119697 240
rect 120239 -480 120295 240
rect 120837 -480 120893 240
rect 121435 -480 121491 240
rect 122033 -480 122089 240
rect 122585 -480 122641 240
rect 123183 -480 123239 240
rect 123781 -480 123837 240
rect 124379 -480 124435 240
rect 124977 -480 125033 240
rect 125575 -480 125631 240
rect 126173 -480 126229 240
rect 126725 -480 126781 240
rect 127323 -480 127379 240
rect 127921 -480 127977 240
rect 128519 -480 128575 240
rect 129117 -480 129173 240
rect 129715 -480 129771 240
rect 130313 -480 130369 240
rect 130865 -480 130921 240
rect 131463 -480 131519 240
rect 132061 -480 132117 240
rect 132659 -480 132715 240
rect 133257 -480 133313 240
rect 133855 -480 133911 240
rect 134407 -480 134463 240
rect 135005 -480 135061 240
rect 135603 -480 135659 240
rect 136201 -480 136257 240
rect 136799 -480 136855 240
rect 137397 -480 137453 240
rect 137995 -480 138051 240
rect 138547 -480 138603 240
rect 139145 -480 139201 240
rect 139743 -480 139799 240
rect 140341 -480 140397 240
rect 140939 -480 140995 240
rect 141537 -480 141593 240
rect 142135 -480 142191 240
rect 142687 -480 142743 240
rect 143285 -480 143341 240
rect 143883 -480 143939 240
rect 144481 -480 144537 240
rect 145079 -480 145135 240
rect 145677 -480 145733 240
rect 146275 -480 146331 240
rect 146827 -480 146883 240
rect 147425 -480 147481 240
rect 148023 -480 148079 240
rect 148621 -480 148677 240
rect 149219 -480 149275 240
rect 149817 -480 149873 240
rect 150369 -480 150425 240
rect 150967 -480 151023 240
rect 151565 -480 151621 240
rect 152163 -480 152219 240
rect 152761 -480 152817 240
rect 153359 -480 153415 240
rect 153957 -480 154013 240
rect 154509 -480 154565 240
rect 155107 -480 155163 240
rect 155705 -480 155761 240
rect 156303 -480 156359 240
rect 156901 -480 156957 240
rect 157499 -480 157555 240
rect 158097 -480 158153 240
rect 158649 -480 158705 240
rect 159247 -480 159303 240
rect 159845 -480 159901 240
rect 160443 -480 160499 240
rect 161041 -480 161097 240
rect 161639 -480 161695 240
rect 162191 -480 162247 240
rect 162789 -480 162845 240
rect 163387 -480 163443 240
rect 163985 -480 164041 240
rect 164583 -480 164639 240
rect 165181 -480 165237 240
rect 165779 -480 165835 240
rect 166331 -480 166387 240
rect 166929 -480 166985 240
rect 167527 -480 167583 240
rect 168125 -480 168181 240
rect 168723 -480 168779 240
rect 169321 -480 169377 240
rect 169919 -480 169975 240
rect 170471 -480 170527 240
rect 171069 -480 171125 240
rect 171667 -480 171723 240
rect 172265 -480 172321 240
rect 172863 -480 172919 240
rect 173461 -480 173517 240
rect 174013 -480 174069 240
rect 174611 -480 174667 240
rect 175209 -480 175265 240
rect 175807 -480 175863 240
rect 176405 -480 176461 240
rect 177003 -480 177059 240
rect 177601 -480 177657 240
rect 178153 -480 178209 240
rect 178751 -480 178807 240
rect 179349 -480 179405 240
rect 179947 -480 180003 240
rect 180545 -480 180601 240
rect 181143 -480 181199 240
rect 181741 -480 181797 240
rect 182293 -480 182349 240
rect 182891 -480 182947 240
rect 183489 -480 183545 240
rect 184087 -480 184143 240
rect 184685 -480 184741 240
rect 185283 -480 185339 240
rect 185835 -480 185891 240
rect 186433 -480 186489 240
rect 187031 -480 187087 240
rect 187629 -480 187685 240
rect 188227 -480 188283 240
rect 188825 -480 188881 240
rect 189423 -480 189479 240
rect 189975 -480 190031 240
rect 190573 -480 190629 240
rect 191171 -480 191227 240
rect 191769 -480 191825 240
rect 192367 -480 192423 240
rect 192965 -480 193021 240
rect 193563 -480 193619 240
rect 194115 -480 194171 240
rect 194713 -480 194769 240
rect 195311 -480 195367 240
rect 195909 -480 195965 240
rect 196507 -480 196563 240
rect 197105 -480 197161 240
rect 197657 -480 197713 240
rect 198255 -480 198311 240
rect 198853 -480 198909 240
rect 199451 -480 199507 240
rect 200049 -480 200105 240
rect 200647 -480 200703 240
rect 201245 -480 201301 240
rect 201797 -480 201853 240
rect 202395 -480 202451 240
rect 202993 -480 203049 240
rect 203591 -480 203647 240
rect 204189 -480 204245 240
rect 204787 -480 204843 240
rect 205385 -480 205441 240
rect 205937 -480 205993 240
rect 206535 -480 206591 240
rect 207133 -480 207189 240
rect 207731 -480 207787 240
rect 208329 -480 208385 240
rect 208927 -480 208983 240
rect 209479 -480 209535 240
rect 210077 -480 210133 240
rect 210675 -480 210731 240
rect 211273 -480 211329 240
rect 211871 -480 211927 240
rect 212469 -480 212525 240
rect 213067 -480 213123 240
rect 213619 -480 213675 240
rect 214217 -480 214273 240
rect 214815 -480 214871 240
rect 215413 -480 215469 240
rect 216011 -480 216067 240
rect 216609 -480 216665 240
rect 217207 -480 217263 240
rect 217759 -480 217815 240
rect 218357 -480 218413 240
rect 218955 -480 219011 240
rect 219553 -480 219609 240
rect 220151 -480 220207 240
rect 220749 -480 220805 240
rect 221301 -480 221357 240
rect 221899 -480 221955 240
rect 222497 -480 222553 240
rect 223095 -480 223151 240
rect 223693 -480 223749 240
rect 224291 -480 224347 240
rect 224889 -480 224945 240
rect 225441 -480 225497 240
rect 226039 -480 226095 240
rect 226637 -480 226693 240
rect 227235 -480 227291 240
rect 227833 -480 227889 240
rect 228431 -480 228487 240
rect 229029 -480 229085 240
rect 229581 -480 229637 240
rect 230179 -480 230235 240
rect 230777 -480 230833 240
rect 231375 -480 231431 240
rect 231973 -480 232029 240
rect 232571 -480 232627 240
rect 233123 -480 233179 240
rect 233721 -480 233777 240
rect 234319 -480 234375 240
rect 234917 -480 234973 240
rect 235515 -480 235571 240
rect 236113 -480 236169 240
rect 236711 -480 236767 240
rect 237263 -480 237319 240
rect 237861 -480 237917 240
rect 238459 -480 238515 240
rect 239057 -480 239113 240
rect 239655 -480 239711 240
rect 240253 -480 240309 240
rect 240851 -480 240907 240
rect 241403 -480 241459 240
rect 242001 -480 242057 240
rect 242599 -480 242655 240
rect 243197 -480 243253 240
rect 243795 -480 243851 240
rect 244393 -480 244449 240
rect 244945 -480 245001 240
rect 245543 -480 245599 240
rect 246141 -480 246197 240
rect 246739 -480 246795 240
rect 247337 -480 247393 240
rect 247935 -480 247991 240
rect 248533 -480 248589 240
rect 249085 -480 249141 240
rect 249683 -480 249739 240
rect 250281 -480 250337 240
rect 250879 -480 250935 240
rect 251477 -480 251533 240
rect 252075 -480 252131 240
rect 252673 -480 252729 240
rect 253225 -480 253281 240
rect 253823 -480 253879 240
rect 254421 -480 254477 240
rect 255019 -480 255075 240
rect 255617 -480 255673 240
rect 256215 -480 256271 240
rect 256767 -480 256823 240
rect 257365 -480 257421 240
rect 257963 -480 258019 240
rect 258561 -480 258617 240
rect 259159 -480 259215 240
rect 259757 -480 259813 240
rect 260355 -480 260411 240
rect 260907 -480 260963 240
rect 261505 -480 261561 240
rect 262103 -480 262159 240
rect 262701 -480 262757 240
rect 263299 -480 263355 240
rect 263897 -480 263953 240
rect 264495 -480 264551 240
rect 265047 -480 265103 240
rect 265645 -480 265701 240
rect 266243 -480 266299 240
rect 266841 -480 266897 240
rect 267439 -480 267495 240
rect 268037 -480 268093 240
rect 268589 -480 268645 240
rect 269187 -480 269243 240
rect 269785 -480 269841 240
rect 270383 -480 270439 240
rect 270981 -480 271037 240
rect 271579 -480 271635 240
rect 272177 -480 272233 240
rect 272729 -480 272785 240
rect 273327 -480 273383 240
rect 273925 -480 273981 240
rect 274523 -480 274579 240
rect 275121 -480 275177 240
rect 275719 -480 275775 240
rect 276317 -480 276373 240
rect 276869 -480 276925 240
rect 277467 -480 277523 240
rect 278065 -480 278121 240
rect 278663 -480 278719 240
rect 279261 -480 279317 240
rect 279859 -480 279915 240
rect 280411 -480 280467 240
rect 281009 -480 281065 240
rect 281607 -480 281663 240
rect 282205 -480 282261 240
rect 282803 -480 282859 240
rect 283401 -480 283457 240
rect 283999 -480 284055 240
rect 284551 -480 284607 240
rect 285149 -480 285205 240
rect 285747 -480 285803 240
rect 286345 -480 286401 240
rect 286943 -480 286999 240
rect 287541 -480 287597 240
rect 288139 -480 288195 240
rect 288691 -480 288747 240
rect 289289 -480 289345 240
rect 289887 -480 289943 240
rect 290485 -480 290541 240
rect 291083 -480 291139 240
rect 291681 -480 291737 240
<< obsm2 >>
rect 286 351732 4015 351760
rect 4127 351732 12111 351760
rect 12223 351732 20207 351760
rect 20319 351732 28349 351760
rect 28461 351732 36445 351760
rect 36557 351732 44541 351760
rect 44653 351732 52683 351760
rect 52795 351732 60779 351760
rect 60891 351732 68875 351760
rect 68987 351732 77017 351760
rect 77129 351732 85113 351760
rect 85225 351732 93209 351760
rect 93321 351732 101351 351760
rect 101463 351732 109447 351760
rect 109559 351732 117543 351760
rect 117655 351732 125685 351760
rect 125797 351732 133781 351760
rect 133893 351732 141877 351760
rect 141989 351732 150019 351760
rect 150131 351732 158115 351760
rect 158227 351732 166211 351760
rect 166323 351732 174353 351760
rect 174465 351732 182449 351760
rect 182561 351732 190545 351760
rect 190657 351732 198687 351760
rect 198799 351732 206783 351760
rect 206895 351732 214879 351760
rect 214991 351732 223021 351760
rect 223133 351732 231117 351760
rect 231229 351732 239213 351760
rect 239325 351732 247355 351760
rect 247467 351732 255451 351760
rect 255563 351732 263547 351760
rect 263659 351732 271689 351760
rect 271801 351732 279785 351760
rect 279897 351732 287881 351760
rect 287993 351732 291814 351760
rect 286 268 291814 351732
rect 355 1 795 268
rect 907 1 1393 268
rect 1505 1 1991 268
rect 2103 1 2589 268
rect 2701 1 3187 268
rect 3299 1 3785 268
rect 3897 1 4337 268
rect 4449 1 4935 268
rect 5047 1 5533 268
rect 5645 1 6131 268
rect 6243 1 6729 268
rect 6841 1 7327 268
rect 7439 1 7925 268
rect 8037 1 8477 268
rect 8589 1 9075 268
rect 9187 1 9673 268
rect 9785 1 10271 268
rect 10383 1 10869 268
rect 10981 1 11467 268
rect 11579 1 12065 268
rect 12177 1 12617 268
rect 12729 1 13215 268
rect 13327 1 13813 268
rect 13925 1 14411 268
rect 14523 1 15009 268
rect 15121 1 15607 268
rect 15719 1 16159 268
rect 16271 1 16757 268
rect 16869 1 17355 268
rect 17467 1 17953 268
rect 18065 1 18551 268
rect 18663 1 19149 268
rect 19261 1 19747 268
rect 19859 1 20299 268
rect 20411 1 20897 268
rect 21009 1 21495 268
rect 21607 1 22093 268
rect 22205 1 22691 268
rect 22803 1 23289 268
rect 23401 1 23887 268
rect 23999 1 24439 268
rect 24551 1 25037 268
rect 25149 1 25635 268
rect 25747 1 26233 268
rect 26345 1 26831 268
rect 26943 1 27429 268
rect 27541 1 27981 268
rect 28093 1 28579 268
rect 28691 1 29177 268
rect 29289 1 29775 268
rect 29887 1 30373 268
rect 30485 1 30971 268
rect 31083 1 31569 268
rect 31681 1 32121 268
rect 32233 1 32719 268
rect 32831 1 33317 268
rect 33429 1 33915 268
rect 34027 1 34513 268
rect 34625 1 35111 268
rect 35223 1 35709 268
rect 35821 1 36261 268
rect 36373 1 36859 268
rect 36971 1 37457 268
rect 37569 1 38055 268
rect 38167 1 38653 268
rect 38765 1 39251 268
rect 39363 1 39803 268
rect 39915 1 40401 268
rect 40513 1 40999 268
rect 41111 1 41597 268
rect 41709 1 42195 268
rect 42307 1 42793 268
rect 42905 1 43391 268
rect 43503 1 43943 268
rect 44055 1 44541 268
rect 44653 1 45139 268
rect 45251 1 45737 268
rect 45849 1 46335 268
rect 46447 1 46933 268
rect 47045 1 47531 268
rect 47643 1 48083 268
rect 48195 1 48681 268
rect 48793 1 49279 268
rect 49391 1 49877 268
rect 49989 1 50475 268
rect 50587 1 51073 268
rect 51185 1 51625 268
rect 51737 1 52223 268
rect 52335 1 52821 268
rect 52933 1 53419 268
rect 53531 1 54017 268
rect 54129 1 54615 268
rect 54727 1 55213 268
rect 55325 1 55765 268
rect 55877 1 56363 268
rect 56475 1 56961 268
rect 57073 1 57559 268
rect 57671 1 58157 268
rect 58269 1 58755 268
rect 58867 1 59353 268
rect 59465 1 59905 268
rect 60017 1 60503 268
rect 60615 1 61101 268
rect 61213 1 61699 268
rect 61811 1 62297 268
rect 62409 1 62895 268
rect 63007 1 63447 268
rect 63559 1 64045 268
rect 64157 1 64643 268
rect 64755 1 65241 268
rect 65353 1 65839 268
rect 65951 1 66437 268
rect 66549 1 67035 268
rect 67147 1 67587 268
rect 67699 1 68185 268
rect 68297 1 68783 268
rect 68895 1 69381 268
rect 69493 1 69979 268
rect 70091 1 70577 268
rect 70689 1 71175 268
rect 71287 1 71727 268
rect 71839 1 72325 268
rect 72437 1 72923 268
rect 73035 1 73521 268
rect 73633 1 74119 268
rect 74231 1 74717 268
rect 74829 1 75269 268
rect 75381 1 75867 268
rect 75979 1 76465 268
rect 76577 1 77063 268
rect 77175 1 77661 268
rect 77773 1 78259 268
rect 78371 1 78857 268
rect 78969 1 79409 268
rect 79521 1 80007 268
rect 80119 1 80605 268
rect 80717 1 81203 268
rect 81315 1 81801 268
rect 81913 1 82399 268
rect 82511 1 82997 268
rect 83109 1 83549 268
rect 83661 1 84147 268
rect 84259 1 84745 268
rect 84857 1 85343 268
rect 85455 1 85941 268
rect 86053 1 86539 268
rect 86651 1 87091 268
rect 87203 1 87689 268
rect 87801 1 88287 268
rect 88399 1 88885 268
rect 88997 1 89483 268
rect 89595 1 90081 268
rect 90193 1 90679 268
rect 90791 1 91231 268
rect 91343 1 91829 268
rect 91941 1 92427 268
rect 92539 1 93025 268
rect 93137 1 93623 268
rect 93735 1 94221 268
rect 94333 1 94819 268
rect 94931 1 95371 268
rect 95483 1 95969 268
rect 96081 1 96567 268
rect 96679 1 97165 268
rect 97277 1 97763 268
rect 97875 1 98361 268
rect 98473 1 98913 268
rect 99025 1 99511 268
rect 99623 1 100109 268
rect 100221 1 100707 268
rect 100819 1 101305 268
rect 101417 1 101903 268
rect 102015 1 102501 268
rect 102613 1 103053 268
rect 103165 1 103651 268
rect 103763 1 104249 268
rect 104361 1 104847 268
rect 104959 1 105445 268
rect 105557 1 106043 268
rect 106155 1 106641 268
rect 106753 1 107193 268
rect 107305 1 107791 268
rect 107903 1 108389 268
rect 108501 1 108987 268
rect 109099 1 109585 268
rect 109697 1 110183 268
rect 110295 1 110735 268
rect 110847 1 111333 268
rect 111445 1 111931 268
rect 112043 1 112529 268
rect 112641 1 113127 268
rect 113239 1 113725 268
rect 113837 1 114323 268
rect 114435 1 114875 268
rect 114987 1 115473 268
rect 115585 1 116071 268
rect 116183 1 116669 268
rect 116781 1 117267 268
rect 117379 1 117865 268
rect 117977 1 118463 268
rect 118575 1 119015 268
rect 119127 1 119613 268
rect 119725 1 120211 268
rect 120323 1 120809 268
rect 120921 1 121407 268
rect 121519 1 122005 268
rect 122117 1 122557 268
rect 122669 1 123155 268
rect 123267 1 123753 268
rect 123865 1 124351 268
rect 124463 1 124949 268
rect 125061 1 125547 268
rect 125659 1 126145 268
rect 126257 1 126697 268
rect 126809 1 127295 268
rect 127407 1 127893 268
rect 128005 1 128491 268
rect 128603 1 129089 268
rect 129201 1 129687 268
rect 129799 1 130285 268
rect 130397 1 130837 268
rect 130949 1 131435 268
rect 131547 1 132033 268
rect 132145 1 132631 268
rect 132743 1 133229 268
rect 133341 1 133827 268
rect 133939 1 134379 268
rect 134491 1 134977 268
rect 135089 1 135575 268
rect 135687 1 136173 268
rect 136285 1 136771 268
rect 136883 1 137369 268
rect 137481 1 137967 268
rect 138079 1 138519 268
rect 138631 1 139117 268
rect 139229 1 139715 268
rect 139827 1 140313 268
rect 140425 1 140911 268
rect 141023 1 141509 268
rect 141621 1 142107 268
rect 142219 1 142659 268
rect 142771 1 143257 268
rect 143369 1 143855 268
rect 143967 1 144453 268
rect 144565 1 145051 268
rect 145163 1 145649 268
rect 145761 1 146247 268
rect 146359 1 146799 268
rect 146911 1 147397 268
rect 147509 1 147995 268
rect 148107 1 148593 268
rect 148705 1 149191 268
rect 149303 1 149789 268
rect 149901 1 150341 268
rect 150453 1 150939 268
rect 151051 1 151537 268
rect 151649 1 152135 268
rect 152247 1 152733 268
rect 152845 1 153331 268
rect 153443 1 153929 268
rect 154041 1 154481 268
rect 154593 1 155079 268
rect 155191 1 155677 268
rect 155789 1 156275 268
rect 156387 1 156873 268
rect 156985 1 157471 268
rect 157583 1 158069 268
rect 158181 1 158621 268
rect 158733 1 159219 268
rect 159331 1 159817 268
rect 159929 1 160415 268
rect 160527 1 161013 268
rect 161125 1 161611 268
rect 161723 1 162163 268
rect 162275 1 162761 268
rect 162873 1 163359 268
rect 163471 1 163957 268
rect 164069 1 164555 268
rect 164667 1 165153 268
rect 165265 1 165751 268
rect 165863 1 166303 268
rect 166415 1 166901 268
rect 167013 1 167499 268
rect 167611 1 168097 268
rect 168209 1 168695 268
rect 168807 1 169293 268
rect 169405 1 169891 268
rect 170003 1 170443 268
rect 170555 1 171041 268
rect 171153 1 171639 268
rect 171751 1 172237 268
rect 172349 1 172835 268
rect 172947 1 173433 268
rect 173545 1 173985 268
rect 174097 1 174583 268
rect 174695 1 175181 268
rect 175293 1 175779 268
rect 175891 1 176377 268
rect 176489 1 176975 268
rect 177087 1 177573 268
rect 177685 1 178125 268
rect 178237 1 178723 268
rect 178835 1 179321 268
rect 179433 1 179919 268
rect 180031 1 180517 268
rect 180629 1 181115 268
rect 181227 1 181713 268
rect 181825 1 182265 268
rect 182377 1 182863 268
rect 182975 1 183461 268
rect 183573 1 184059 268
rect 184171 1 184657 268
rect 184769 1 185255 268
rect 185367 1 185807 268
rect 185919 1 186405 268
rect 186517 1 187003 268
rect 187115 1 187601 268
rect 187713 1 188199 268
rect 188311 1 188797 268
rect 188909 1 189395 268
rect 189507 1 189947 268
rect 190059 1 190545 268
rect 190657 1 191143 268
rect 191255 1 191741 268
rect 191853 1 192339 268
rect 192451 1 192937 268
rect 193049 1 193535 268
rect 193647 1 194087 268
rect 194199 1 194685 268
rect 194797 1 195283 268
rect 195395 1 195881 268
rect 195993 1 196479 268
rect 196591 1 197077 268
rect 197189 1 197629 268
rect 197741 1 198227 268
rect 198339 1 198825 268
rect 198937 1 199423 268
rect 199535 1 200021 268
rect 200133 1 200619 268
rect 200731 1 201217 268
rect 201329 1 201769 268
rect 201881 1 202367 268
rect 202479 1 202965 268
rect 203077 1 203563 268
rect 203675 1 204161 268
rect 204273 1 204759 268
rect 204871 1 205357 268
rect 205469 1 205909 268
rect 206021 1 206507 268
rect 206619 1 207105 268
rect 207217 1 207703 268
rect 207815 1 208301 268
rect 208413 1 208899 268
rect 209011 1 209451 268
rect 209563 1 210049 268
rect 210161 1 210647 268
rect 210759 1 211245 268
rect 211357 1 211843 268
rect 211955 1 212441 268
rect 212553 1 213039 268
rect 213151 1 213591 268
rect 213703 1 214189 268
rect 214301 1 214787 268
rect 214899 1 215385 268
rect 215497 1 215983 268
rect 216095 1 216581 268
rect 216693 1 217179 268
rect 217291 1 217731 268
rect 217843 1 218329 268
rect 218441 1 218927 268
rect 219039 1 219525 268
rect 219637 1 220123 268
rect 220235 1 220721 268
rect 220833 1 221273 268
rect 221385 1 221871 268
rect 221983 1 222469 268
rect 222581 1 223067 268
rect 223179 1 223665 268
rect 223777 1 224263 268
rect 224375 1 224861 268
rect 224973 1 225413 268
rect 225525 1 226011 268
rect 226123 1 226609 268
rect 226721 1 227207 268
rect 227319 1 227805 268
rect 227917 1 228403 268
rect 228515 1 229001 268
rect 229113 1 229553 268
rect 229665 1 230151 268
rect 230263 1 230749 268
rect 230861 1 231347 268
rect 231459 1 231945 268
rect 232057 1 232543 268
rect 232655 1 233095 268
rect 233207 1 233693 268
rect 233805 1 234291 268
rect 234403 1 234889 268
rect 235001 1 235487 268
rect 235599 1 236085 268
rect 236197 1 236683 268
rect 236795 1 237235 268
rect 237347 1 237833 268
rect 237945 1 238431 268
rect 238543 1 239029 268
rect 239141 1 239627 268
rect 239739 1 240225 268
rect 240337 1 240823 268
rect 240935 1 241375 268
rect 241487 1 241973 268
rect 242085 1 242571 268
rect 242683 1 243169 268
rect 243281 1 243767 268
rect 243879 1 244365 268
rect 244477 1 244917 268
rect 245029 1 245515 268
rect 245627 1 246113 268
rect 246225 1 246711 268
rect 246823 1 247309 268
rect 247421 1 247907 268
rect 248019 1 248505 268
rect 248617 1 249057 268
rect 249169 1 249655 268
rect 249767 1 250253 268
rect 250365 1 250851 268
rect 250963 1 251449 268
rect 251561 1 252047 268
rect 252159 1 252645 268
rect 252757 1 253197 268
rect 253309 1 253795 268
rect 253907 1 254393 268
rect 254505 1 254991 268
rect 255103 1 255589 268
rect 255701 1 256187 268
rect 256299 1 256739 268
rect 256851 1 257337 268
rect 257449 1 257935 268
rect 258047 1 258533 268
rect 258645 1 259131 268
rect 259243 1 259729 268
rect 259841 1 260327 268
rect 260439 1 260879 268
rect 260991 1 261477 268
rect 261589 1 262075 268
rect 262187 1 262673 268
rect 262785 1 263271 268
rect 263383 1 263869 268
rect 263981 1 264467 268
rect 264579 1 265019 268
rect 265131 1 265617 268
rect 265729 1 266215 268
rect 266327 1 266813 268
rect 266925 1 267411 268
rect 267523 1 268009 268
rect 268121 1 268561 268
rect 268673 1 269159 268
rect 269271 1 269757 268
rect 269869 1 270355 268
rect 270467 1 270953 268
rect 271065 1 271551 268
rect 271663 1 272149 268
rect 272261 1 272701 268
rect 272813 1 273299 268
rect 273411 1 273897 268
rect 274009 1 274495 268
rect 274607 1 275093 268
rect 275205 1 275691 268
rect 275803 1 276289 268
rect 276401 1 276841 268
rect 276953 1 277439 268
rect 277551 1 278037 268
rect 278149 1 278635 268
rect 278747 1 279233 268
rect 279345 1 279831 268
rect 279943 1 280383 268
rect 280495 1 280981 268
rect 281093 1 281579 268
rect 281691 1 282177 268
rect 282289 1 282775 268
rect 282887 1 283373 268
rect 283485 1 283971 268
rect 284083 1 284523 268
rect 284635 1 285121 268
rect 285233 1 285719 268
rect 285831 1 286317 268
rect 286429 1 286915 268
rect 287027 1 287513 268
rect 287625 1 288111 268
rect 288223 1 288663 268
rect 288775 1 289261 268
rect 289373 1 289859 268
rect 289971 1 290457 268
rect 290569 1 291055 268
rect 291167 1 291653 268
rect 291765 1 291814 268
<< metal3 >>
rect -480 348610 240 348730
rect 291760 348542 292480 348662
rect -480 342082 240 342202
rect 291760 341878 292480 341998
rect -480 335554 240 335674
rect 291760 335282 292480 335402
rect -480 329026 240 329146
rect 291760 328618 292480 328738
rect -480 322498 240 322618
rect 291760 321954 292480 322074
rect -480 315970 240 316090
rect 291760 315358 292480 315478
rect -480 309510 240 309630
rect 291760 308694 292480 308814
rect -480 302982 240 303102
rect 291760 302030 292480 302150
rect -480 296454 240 296574
rect 291760 295434 292480 295554
rect -480 289926 240 290046
rect 291760 288770 292480 288890
rect -480 283398 240 283518
rect 291760 282106 292480 282226
rect -480 276870 240 276990
rect 291760 275510 292480 275630
rect -480 270342 240 270462
rect 291760 268846 292480 268966
rect -480 263882 240 264002
rect 291760 262182 292480 262302
rect -480 257354 240 257474
rect 291760 255586 292480 255706
rect -480 250826 240 250946
rect 291760 248922 292480 249042
rect -480 244298 240 244418
rect 291760 242258 292480 242378
rect -480 237770 240 237890
rect 291760 235662 292480 235782
rect -480 231242 240 231362
rect 291760 228998 292480 229118
rect -480 224714 240 224834
rect 291760 222334 292480 222454
rect -480 218254 240 218374
rect 291760 215738 292480 215858
rect -480 211726 240 211846
rect 291760 209074 292480 209194
rect -480 205198 240 205318
rect 291760 202410 292480 202530
rect -480 198670 240 198790
rect 291760 195814 292480 195934
rect -480 192142 240 192262
rect 291760 189150 292480 189270
rect -480 185614 240 185734
rect 291760 182486 292480 182606
rect -480 179154 240 179274
rect 291760 175890 292480 176010
rect -480 172626 240 172746
rect 291760 169226 292480 169346
rect -480 166098 240 166218
rect 291760 162562 292480 162682
rect -480 159570 240 159690
rect 291760 155966 292480 156086
rect -480 153042 240 153162
rect 291760 149302 292480 149422
rect -480 146514 240 146634
rect 291760 142638 292480 142758
rect -480 139986 240 140106
rect 291760 136042 292480 136162
rect -480 133526 240 133646
rect 291760 129378 292480 129498
rect -480 126998 240 127118
rect 291760 122714 292480 122834
rect -480 120470 240 120590
rect 291760 116118 292480 116238
rect -480 113942 240 114062
rect 291760 109454 292480 109574
rect -480 107414 240 107534
rect 291760 102790 292480 102910
rect -480 100886 240 101006
rect 291760 96194 292480 96314
rect -480 94358 240 94478
rect 291760 89530 292480 89650
rect -480 87898 240 88018
rect 291760 82866 292480 82986
rect -480 81370 240 81490
rect 291760 76270 292480 76390
rect -480 74842 240 74962
rect 291760 69606 292480 69726
rect -480 68314 240 68434
rect 291760 62942 292480 63062
rect -480 61786 240 61906
rect 291760 56346 292480 56466
rect -480 55258 240 55378
rect 291760 49682 292480 49802
rect -480 48730 240 48850
rect 291760 43018 292480 43138
rect -480 42270 240 42390
rect 291760 36422 292480 36542
rect -480 35742 240 35862
rect 291760 29758 292480 29878
rect -480 29214 240 29334
rect 291760 23094 292480 23214
rect -480 22686 240 22806
rect 291760 16498 292480 16618
rect -480 16158 240 16278
rect 291760 9834 292480 9954
rect -480 9630 240 9750
rect -480 3170 240 3290
rect 291760 3238 292480 3358
<< obsm3 >>
rect 240 348770 291793 349004
rect 280 348702 291793 348770
rect 280 348570 291720 348702
rect 240 348502 291720 348570
rect 240 342242 291793 348502
rect 280 342042 291793 342242
rect 240 342038 291793 342042
rect 240 341838 291720 342038
rect 240 335714 291793 341838
rect 280 335514 291793 335714
rect 240 335442 291793 335514
rect 240 335242 291720 335442
rect 240 329186 291793 335242
rect 280 328986 291793 329186
rect 240 328778 291793 328986
rect 240 328578 291720 328778
rect 240 322658 291793 328578
rect 280 322458 291793 322658
rect 240 322114 291793 322458
rect 240 321914 291720 322114
rect 240 316130 291793 321914
rect 280 315930 291793 316130
rect 240 315518 291793 315930
rect 240 315318 291720 315518
rect 240 309670 291793 315318
rect 280 309470 291793 309670
rect 240 308854 291793 309470
rect 240 308654 291720 308854
rect 240 303142 291793 308654
rect 280 302942 291793 303142
rect 240 302190 291793 302942
rect 240 301990 291720 302190
rect 240 296614 291793 301990
rect 280 296414 291793 296614
rect 240 295594 291793 296414
rect 240 295394 291720 295594
rect 240 290086 291793 295394
rect 280 289886 291793 290086
rect 240 288930 291793 289886
rect 240 288730 291720 288930
rect 240 283558 291793 288730
rect 280 283358 291793 283558
rect 240 282266 291793 283358
rect 240 282066 291720 282266
rect 240 277030 291793 282066
rect 280 276830 291793 277030
rect 240 275670 291793 276830
rect 240 275470 291720 275670
rect 240 270502 291793 275470
rect 280 270302 291793 270502
rect 240 269006 291793 270302
rect 240 268806 291720 269006
rect 240 264042 291793 268806
rect 280 263842 291793 264042
rect 240 262342 291793 263842
rect 240 262142 291720 262342
rect 240 257514 291793 262142
rect 280 257314 291793 257514
rect 240 255746 291793 257314
rect 240 255546 291720 255746
rect 240 250986 291793 255546
rect 280 250786 291793 250986
rect 240 249082 291793 250786
rect 240 248882 291720 249082
rect 240 244458 291793 248882
rect 280 244258 291793 244458
rect 240 242418 291793 244258
rect 240 242218 291720 242418
rect 240 237930 291793 242218
rect 280 237730 291793 237930
rect 240 235822 291793 237730
rect 240 235622 291720 235822
rect 240 231402 291793 235622
rect 280 231202 291793 231402
rect 240 229158 291793 231202
rect 240 228958 291720 229158
rect 240 224874 291793 228958
rect 280 224674 291793 224874
rect 240 222494 291793 224674
rect 240 222294 291720 222494
rect 240 218414 291793 222294
rect 280 218214 291793 218414
rect 240 215898 291793 218214
rect 240 215698 291720 215898
rect 240 211886 291793 215698
rect 280 211686 291793 211886
rect 240 209234 291793 211686
rect 240 209034 291720 209234
rect 240 205358 291793 209034
rect 280 205158 291793 205358
rect 240 202570 291793 205158
rect 240 202370 291720 202570
rect 240 198830 291793 202370
rect 280 198630 291793 198830
rect 240 195974 291793 198630
rect 240 195774 291720 195974
rect 240 192302 291793 195774
rect 280 192102 291793 192302
rect 240 189310 291793 192102
rect 240 189110 291720 189310
rect 240 185774 291793 189110
rect 280 185574 291793 185774
rect 240 182646 291793 185574
rect 240 182446 291720 182646
rect 240 179314 291793 182446
rect 280 179114 291793 179314
rect 240 176050 291793 179114
rect 240 175850 291720 176050
rect 240 172786 291793 175850
rect 280 172586 291793 172786
rect 240 169386 291793 172586
rect 240 169186 291720 169386
rect 240 166258 291793 169186
rect 280 166058 291793 166258
rect 240 162722 291793 166058
rect 240 162522 291720 162722
rect 240 159730 291793 162522
rect 280 159530 291793 159730
rect 240 156126 291793 159530
rect 240 155926 291720 156126
rect 240 153202 291793 155926
rect 280 153002 291793 153202
rect 240 149462 291793 153002
rect 240 149262 291720 149462
rect 240 146674 291793 149262
rect 280 146474 291793 146674
rect 240 142798 291793 146474
rect 240 142598 291720 142798
rect 240 140146 291793 142598
rect 280 139946 291793 140146
rect 240 136202 291793 139946
rect 240 136002 291720 136202
rect 240 133686 291793 136002
rect 280 133486 291793 133686
rect 240 129538 291793 133486
rect 240 129338 291720 129538
rect 240 127158 291793 129338
rect 280 126958 291793 127158
rect 240 122874 291793 126958
rect 240 122674 291720 122874
rect 240 120630 291793 122674
rect 280 120430 291793 120630
rect 240 116278 291793 120430
rect 240 116078 291720 116278
rect 240 114102 291793 116078
rect 280 113902 291793 114102
rect 240 109614 291793 113902
rect 240 109414 291720 109614
rect 240 107574 291793 109414
rect 280 107374 291793 107574
rect 240 102950 291793 107374
rect 240 102750 291720 102950
rect 240 101046 291793 102750
rect 280 100846 291793 101046
rect 240 96354 291793 100846
rect 240 96154 291720 96354
rect 240 94518 291793 96154
rect 280 94318 291793 94518
rect 240 89690 291793 94318
rect 240 89490 291720 89690
rect 240 88058 291793 89490
rect 280 87858 291793 88058
rect 240 83026 291793 87858
rect 240 82826 291720 83026
rect 240 81530 291793 82826
rect 280 81330 291793 81530
rect 240 76430 291793 81330
rect 240 76230 291720 76430
rect 240 75002 291793 76230
rect 280 74802 291793 75002
rect 240 69766 291793 74802
rect 240 69566 291720 69766
rect 240 68474 291793 69566
rect 280 68274 291793 68474
rect 240 63102 291793 68274
rect 240 62902 291720 63102
rect 240 61946 291793 62902
rect 280 61746 291793 61946
rect 240 56506 291793 61746
rect 240 56306 291720 56506
rect 240 55418 291793 56306
rect 280 55218 291793 55418
rect 240 49842 291793 55218
rect 240 49642 291720 49842
rect 240 48890 291793 49642
rect 280 48690 291793 48890
rect 240 43178 291793 48690
rect 240 42978 291720 43178
rect 240 42430 291793 42978
rect 280 42230 291793 42430
rect 240 36582 291793 42230
rect 240 36382 291720 36582
rect 240 35902 291793 36382
rect 280 35702 291793 35902
rect 240 29918 291793 35702
rect 240 29718 291720 29918
rect 240 29374 291793 29718
rect 280 29174 291793 29374
rect 240 23254 291793 29174
rect 240 23054 291720 23254
rect 240 22846 291793 23054
rect 280 22646 291793 22846
rect 240 16658 291793 22646
rect 240 16458 291720 16658
rect 240 16318 291793 16458
rect 280 16118 291793 16318
rect 240 9994 291793 16118
rect 240 9794 291720 9994
rect 240 9790 291793 9794
rect 280 9590 291793 9790
rect 240 3398 291793 9590
rect 240 3330 291720 3398
rect 280 3198 291720 3330
rect 280 3130 291793 3198
rect 240 2000 291793 3130
<< metal4 >>
rect -4363 -3827 -4053 355795
rect -3883 -3347 -3573 355315
rect -3403 -2867 -3093 354835
rect -2923 -2387 -2613 354355
rect -2443 -1907 -2133 353875
rect -1963 -1427 -1653 353395
rect -1483 -947 -1173 352915
rect -1003 -467 -693 352435
rect 897 350004 1207 352915
rect 2757 350004 3067 353875
rect 4617 350004 4927 354835
rect 6477 350004 6787 355795
rect 9897 350004 10207 352915
rect 11757 350004 12067 353875
rect 13617 350004 13927 354835
rect 15477 350004 15787 355795
rect 18897 350004 19207 352915
rect 20757 350004 21067 353875
rect 22617 350004 22927 354835
rect 24477 350004 24787 355795
rect 27897 350004 28207 352915
rect 29757 350004 30067 353875
rect 31617 350004 31927 354835
rect 33477 350004 33787 355795
rect 36897 350004 37207 352915
rect 38757 350004 39067 353875
rect 40617 350004 40927 354835
rect 42477 350004 42787 355795
rect 45897 350004 46207 352915
rect 47757 350004 48067 353875
rect 49617 350004 49927 354835
rect 51477 350004 51787 355795
rect 54897 350004 55207 352915
rect 56757 350004 57067 353875
rect 58617 350004 58927 354835
rect 60477 350004 60787 355795
rect 63897 350004 64207 352915
rect 65757 350004 66067 353875
rect 67617 350004 67927 354835
rect 69477 350004 69787 355795
rect 72897 350004 73207 352915
rect 74757 350004 75067 353875
rect 76617 350004 76927 354835
rect 78477 350004 78787 355795
rect 81897 350004 82207 352915
rect 83757 350004 84067 353875
rect 85617 350004 85927 354835
rect 87477 350004 87787 355795
rect 90897 350004 91207 352915
rect 92757 350004 93067 353875
rect 94617 350004 94927 354835
rect 96477 350004 96787 355795
rect 99897 350004 100207 352915
rect 101757 350004 102067 353875
rect 103617 350004 103927 354835
rect 105477 350004 105787 355795
rect 108897 350004 109207 352915
rect 110757 350004 111067 353875
rect 112617 350004 112927 354835
rect 114477 350004 114787 355795
rect 117897 350004 118207 352915
rect 119757 350004 120067 353875
rect 121617 350004 121927 354835
rect 123477 350004 123787 355795
rect 126897 350004 127207 352915
rect 128757 350004 129067 353875
rect 130617 350004 130927 354835
rect 132477 350004 132787 355795
rect 135897 350004 136207 352915
rect 137757 350004 138067 353875
rect 139617 350004 139927 354835
rect 141477 350004 141787 355795
rect 144897 350004 145207 352915
rect 146757 350004 147067 353875
rect 148617 350004 148927 354835
rect 150477 350004 150787 355795
rect 153897 350004 154207 352915
rect 155757 350004 156067 353875
rect 157617 350004 157927 354835
rect 159477 350004 159787 355795
rect 162897 350004 163207 352915
rect 164757 350004 165067 353875
rect 166617 350004 166927 354835
rect 168477 350004 168787 355795
rect 171897 350004 172207 352915
rect 173757 350004 174067 353875
rect 175617 350004 175927 354835
rect 177477 350004 177787 355795
rect 180897 350004 181207 352915
rect 182757 350004 183067 353875
rect 184617 350004 184927 354835
rect 186477 350004 186787 355795
rect 189897 350004 190207 352915
rect 191757 350004 192067 353875
rect 193617 350004 193927 354835
rect 195477 350004 195787 355795
rect 198897 350004 199207 352915
rect 200757 350004 201067 353875
rect 202617 350004 202927 354835
rect 204477 350004 204787 355795
rect 207897 350004 208207 352915
rect 209757 350004 210067 353875
rect 211617 350004 211927 354835
rect 213477 350004 213787 355795
rect 216897 350004 217207 352915
rect 218757 350004 219067 353875
rect 220617 350004 220927 354835
rect 222477 350004 222787 355795
rect 225897 350004 226207 352915
rect 227757 350004 228067 353875
rect 229617 350004 229927 354835
rect 231477 350004 231787 355795
rect 234897 350004 235207 352915
rect 236757 350004 237067 353875
rect 238617 350004 238927 354835
rect 240477 350004 240787 355795
rect 243897 350004 244207 352915
rect 245757 350004 246067 353875
rect 247617 350004 247927 354835
rect 249477 350004 249787 355795
rect 252897 350004 253207 352915
rect 254757 350004 255067 353875
rect 256617 350004 256927 354835
rect 258477 350004 258787 355795
rect 261897 350004 262207 352915
rect 263757 350004 264067 353875
rect 265617 350004 265927 354835
rect 267477 350004 267787 355795
rect 270897 350004 271207 352915
rect 272757 350004 273067 353875
rect 274617 350004 274927 354835
rect 276477 350004 276787 355795
rect 279897 350004 280207 352915
rect 281757 350004 282067 353875
rect 283617 350004 283927 354835
rect 285477 350004 285787 355795
rect 288897 350004 289207 352915
rect 897 -947 1207 1000
rect 2757 -1907 3067 1000
rect 4617 -2867 4927 1000
rect 6477 -3827 6787 1000
rect 9897 -947 10207 1000
rect 11757 -1907 12067 1000
rect 13617 -2867 13927 1000
rect 15477 -3827 15787 1000
rect 18897 -947 19207 1000
rect 20757 -1907 21067 1000
rect 22617 -2867 22927 1000
rect 24477 -3827 24787 1000
rect 27897 -947 28207 1000
rect 29757 -1907 30067 1000
rect 31617 -2867 31927 1000
rect 33477 -3827 33787 1000
rect 36897 -947 37207 1000
rect 38757 -1907 39067 1000
rect 40617 -2867 40927 1000
rect 42477 -3827 42787 1000
rect 45897 -947 46207 1000
rect 47757 -1907 48067 1000
rect 49617 -2867 49927 1000
rect 51477 -3827 51787 1000
rect 54897 -947 55207 1000
rect 56757 -1907 57067 1000
rect 58617 -2867 58927 1000
rect 60477 -3827 60787 1000
rect 63897 -947 64207 1000
rect 65757 -1907 66067 1000
rect 67617 -2867 67927 1000
rect 69477 -3827 69787 1000
rect 72897 -947 73207 1000
rect 74757 -1907 75067 1000
rect 76617 -2867 76927 1000
rect 78477 -3827 78787 1000
rect 81897 -947 82207 1000
rect 83757 -1907 84067 1000
rect 85617 -2867 85927 1000
rect 87477 -3827 87787 1000
rect 90897 -947 91207 1000
rect 92757 -1907 93067 1000
rect 94617 -2867 94927 1000
rect 96477 -3827 96787 1000
rect 99897 -947 100207 1000
rect 101757 -1907 102067 1000
rect 103617 -2867 103927 1000
rect 105477 -3827 105787 1000
rect 108897 -947 109207 1000
rect 110757 -1907 111067 1000
rect 112617 -2867 112927 1000
rect 114477 -3827 114787 1000
rect 117897 -947 118207 1000
rect 119757 -1907 120067 1000
rect 121617 -2867 121927 1000
rect 123477 -3827 123787 1000
rect 126897 -947 127207 1000
rect 128757 -1907 129067 1000
rect 130617 -2867 130927 1000
rect 132477 -3827 132787 1000
rect 135897 -947 136207 1000
rect 137757 -1907 138067 1000
rect 139617 -2867 139927 1000
rect 141477 -3827 141787 1000
rect 144897 -947 145207 1000
rect 146757 -1907 147067 1000
rect 148617 -2867 148927 1000
rect 150477 -3827 150787 1000
rect 153897 -947 154207 1000
rect 155757 -1907 156067 1000
rect 157617 -2867 157927 1000
rect 159477 -3827 159787 1000
rect 162897 -947 163207 1000
rect 164757 -1907 165067 1000
rect 166617 -2867 166927 1000
rect 168477 -3827 168787 1000
rect 171897 -947 172207 1000
rect 173757 -1907 174067 1000
rect 175617 -2867 175927 1000
rect 177477 -3827 177787 1000
rect 180897 -947 181207 1000
rect 182757 -1907 183067 1000
rect 184617 -2867 184927 1000
rect 186477 -3827 186787 1000
rect 189897 -947 190207 1000
rect 191757 -1907 192067 1000
rect 193617 -2867 193927 1000
rect 195477 -3827 195787 1000
rect 198897 -947 199207 1000
rect 200757 -1907 201067 1000
rect 202617 -2867 202927 1000
rect 204477 -3827 204787 1000
rect 207897 -947 208207 1000
rect 209757 -1907 210067 1000
rect 211617 -2867 211927 1000
rect 213477 -3827 213787 1000
rect 216897 -947 217207 1000
rect 218757 -1907 219067 1000
rect 220617 -2867 220927 1000
rect 222477 -3827 222787 1000
rect 225897 -947 226207 1000
rect 227757 -1907 228067 1000
rect 229617 -2867 229927 1000
rect 231477 -3827 231787 1000
rect 234897 -947 235207 1000
rect 236757 -1907 237067 1000
rect 238617 -2867 238927 1000
rect 240477 -3827 240787 1000
rect 243897 -947 244207 1000
rect 245757 -1907 246067 1000
rect 247617 -2867 247927 1000
rect 249477 -3827 249787 1000
rect 252897 -947 253207 1000
rect 254757 -1907 255067 1000
rect 256617 -2867 256927 1000
rect 258477 -3827 258787 1000
rect 261897 -947 262207 1000
rect 263757 -1907 264067 1000
rect 265617 -2867 265927 1000
rect 267477 -3827 267787 1000
rect 270897 -947 271207 1000
rect 272757 -1907 273067 1000
rect 274617 -2867 274927 1000
rect 276477 -3827 276787 1000
rect 279897 -947 280207 1000
rect 281757 -1907 282067 1000
rect 283617 -2867 283927 1000
rect 285477 -3827 285787 1000
rect 288897 -947 289207 1000
rect 290757 -1907 291067 353875
rect 292655 -467 292965 352435
rect 293135 -947 293445 352915
rect 293615 -1427 293925 353395
rect 294095 -1907 294405 353875
rect 294575 -2387 294885 354355
rect 295055 -2867 295365 354835
rect 295535 -3347 295845 355315
rect 296015 -3827 296325 355795
<< obsm4 >>
rect 2000 2000 287982 349004
<< metal5 >>
rect -4363 355485 296325 355795
rect -3883 355005 295845 355315
rect -3403 354525 295365 354835
rect -2923 354045 294885 354355
rect -2443 353565 294405 353875
rect -1963 353085 293925 353395
rect -1483 352605 293445 352915
rect -1003 352125 292965 352435
rect -4363 349013 296325 349323
rect -3403 347153 295365 347463
rect -2443 345293 294405 345603
rect -1483 343433 293445 343743
rect -4363 340013 296325 340323
rect -3403 338153 295365 338463
rect -2443 336293 294405 336603
rect -1483 334433 293445 334743
rect -4363 331013 296325 331323
rect -3403 329153 295365 329463
rect -2443 327293 294405 327603
rect -1483 325433 293445 325743
rect -4363 322013 296325 322323
rect -3403 320153 295365 320463
rect -2443 318293 294405 318603
rect -1483 316433 293445 316743
rect -4363 313013 296325 313323
rect -3403 311153 295365 311463
rect -2443 309293 294405 309603
rect -1483 307433 293445 307743
rect -4363 304013 296325 304323
rect -3403 302153 295365 302463
rect -2443 300293 294405 300603
rect -1483 298433 293445 298743
rect -4363 295013 296325 295323
rect -3403 293153 295365 293463
rect -2443 291293 294405 291603
rect -1483 289433 293445 289743
rect -4363 286013 296325 286323
rect -3403 284153 295365 284463
rect -2443 282293 294405 282603
rect -1483 280433 293445 280743
rect -4363 277013 296325 277323
rect -3403 275153 295365 275463
rect -2443 273293 294405 273603
rect -1483 271433 293445 271743
rect -4363 268013 296325 268323
rect -3403 266153 295365 266463
rect -2443 264293 294405 264603
rect -1483 262433 293445 262743
rect -4363 259013 296325 259323
rect -3403 257153 295365 257463
rect -2443 255293 294405 255603
rect -1483 253433 293445 253743
rect -4363 250013 296325 250323
rect -3403 248153 295365 248463
rect -2443 246293 294405 246603
rect -1483 244433 293445 244743
rect -4363 241013 296325 241323
rect -3403 239153 295365 239463
rect -2443 237293 294405 237603
rect -1483 235433 293445 235743
rect -4363 232013 296325 232323
rect -3403 230153 295365 230463
rect -2443 228293 294405 228603
rect -1483 226433 293445 226743
rect -4363 223013 296325 223323
rect -3403 221153 295365 221463
rect -2443 219293 294405 219603
rect -1483 217433 293445 217743
rect -4363 214013 296325 214323
rect -3403 212153 295365 212463
rect -2443 210293 294405 210603
rect -1483 208433 293445 208743
rect -4363 205013 296325 205323
rect -3403 203153 295365 203463
rect -2443 201293 294405 201603
rect -1483 199433 293445 199743
rect -4363 196013 296325 196323
rect -3403 194153 295365 194463
rect -2443 192293 294405 192603
rect -1483 190433 293445 190743
rect -4363 187013 296325 187323
rect -3403 185153 295365 185463
rect -2443 183293 294405 183603
rect -1483 181433 293445 181743
rect -4363 178013 296325 178323
rect -3403 176153 295365 176463
rect -2443 174293 294405 174603
rect -1483 172433 293445 172743
rect -4363 169013 296325 169323
rect -3403 167153 295365 167463
rect -2443 165293 294405 165603
rect -1483 163433 293445 163743
rect -4363 160013 296325 160323
rect -3403 158153 295365 158463
rect -2443 156293 294405 156603
rect -1483 154433 293445 154743
rect -4363 151013 296325 151323
rect -3403 149153 295365 149463
rect -2443 147293 294405 147603
rect -1483 145433 293445 145743
rect -4363 142013 296325 142323
rect -3403 140153 295365 140463
rect -2443 138293 294405 138603
rect -1483 136433 293445 136743
rect -4363 133013 296325 133323
rect -3403 131153 295365 131463
rect -2443 129293 294405 129603
rect -1483 127433 293445 127743
rect -4363 124013 296325 124323
rect -3403 122153 295365 122463
rect -2443 120293 294405 120603
rect -1483 118433 293445 118743
rect -4363 115013 296325 115323
rect -3403 113153 295365 113463
rect -2443 111293 294405 111603
rect -1483 109433 293445 109743
rect -4363 106013 296325 106323
rect -3403 104153 295365 104463
rect -2443 102293 294405 102603
rect -1483 100433 293445 100743
rect -4363 97013 296325 97323
rect -3403 95153 295365 95463
rect -2443 93293 294405 93603
rect -1483 91433 293445 91743
rect -4363 88013 296325 88323
rect -3403 86153 295365 86463
rect -2443 84293 294405 84603
rect -1483 82433 293445 82743
rect -4363 79013 296325 79323
rect -3403 77153 295365 77463
rect -2443 75293 294405 75603
rect -1483 73433 293445 73743
rect -4363 70013 296325 70323
rect -3403 68153 295365 68463
rect -2443 66293 294405 66603
rect -1483 64433 293445 64743
rect -4363 61013 296325 61323
rect -3403 59153 295365 59463
rect -2443 57293 294405 57603
rect -1483 55433 293445 55743
rect -4363 52013 296325 52323
rect -3403 50153 295365 50463
rect -2443 48293 294405 48603
rect -1483 46433 293445 46743
rect -4363 43013 296325 43323
rect -3403 41153 295365 41463
rect -2443 39293 294405 39603
rect -1483 37433 293445 37743
rect -4363 34013 296325 34323
rect -3403 32153 295365 32463
rect -2443 30293 294405 30603
rect -1483 28433 293445 28743
rect -4363 25013 296325 25323
rect -3403 23153 295365 23463
rect -2443 21293 294405 21603
rect -1483 19433 293445 19743
rect -4363 16013 296325 16323
rect -3403 14153 295365 14463
rect -2443 12293 294405 12603
rect -1483 10433 293445 10743
rect -4363 7013 296325 7323
rect -3403 5153 295365 5463
rect -2443 3293 294405 3603
rect -1483 1433 293445 1743
rect -1003 -467 292965 -157
rect -1483 -947 293445 -637
rect -1963 -1427 293925 -1117
rect -2443 -1907 294405 -1597
rect -2923 -2387 294885 -2077
rect -3403 -2867 295365 -2557
rect -3883 -3347 295845 -3037
rect -4363 -3827 296325 -3517
<< obsm5 >>
rect 2000 345763 287982 346874
rect 2000 343903 287982 345133
rect 2000 340483 287982 343273
rect 2000 338623 287982 339853
rect 2000 336763 287982 337993
rect 2000 334903 287982 336133
rect 2000 331483 287982 334273
rect 2000 329623 287982 330853
rect 2000 327763 287982 328993
rect 2000 325903 287982 327133
rect 2000 322483 287982 325273
rect 2000 320623 287982 321853
rect 2000 318763 287982 319993
rect 2000 316903 287982 318133
rect 2000 313483 287982 316273
rect 2000 311623 287982 312853
rect 2000 309763 287982 310993
rect 2000 307903 287982 309133
rect 2000 304483 287982 307273
rect 2000 302623 287982 303853
rect 2000 300763 287982 301993
rect 2000 298903 287982 300133
rect 2000 295483 287982 298273
rect 2000 293623 287982 294853
rect 2000 291763 287982 292993
rect 2000 289903 287982 291133
rect 2000 286483 287982 289273
rect 2000 284623 287982 285853
rect 2000 282763 287982 283993
rect 2000 280903 287982 282133
rect 2000 277483 287982 280273
rect 2000 275623 287982 276853
rect 2000 273763 287982 274993
rect 2000 271903 287982 273133
rect 2000 268483 287982 271273
rect 2000 266623 287982 267853
rect 2000 264763 287982 265993
rect 2000 262903 287982 264133
rect 2000 259483 287982 262273
rect 2000 257623 287982 258853
rect 2000 255763 287982 256993
rect 2000 253903 287982 255133
rect 2000 250483 287982 253273
rect 2000 248623 287982 249853
rect 2000 246763 287982 247993
rect 2000 244903 287982 246133
rect 2000 241483 287982 244273
rect 2000 239623 287982 240853
rect 2000 237763 287982 238993
rect 2000 235903 287982 237133
rect 2000 232483 287982 235273
rect 2000 230623 287982 231853
rect 2000 228763 287982 229993
rect 2000 226903 287982 228133
rect 2000 223483 287982 226273
rect 2000 221623 287982 222853
rect 2000 219763 287982 220993
rect 2000 217903 287982 219133
rect 2000 214483 287982 217273
rect 2000 212623 287982 213853
rect 2000 210763 287982 211993
rect 2000 208903 287982 210133
rect 2000 205483 287982 208273
rect 2000 203623 287982 204853
rect 2000 201763 287982 202993
rect 2000 199903 287982 201133
rect 2000 196483 287982 199273
rect 2000 194623 287982 195853
rect 2000 192763 287982 193993
rect 2000 190903 287982 192133
rect 2000 187483 287982 190273
rect 2000 185623 287982 186853
rect 2000 183763 287982 184993
rect 2000 181903 287982 183133
rect 2000 178483 287982 181273
rect 2000 176623 287982 177853
rect 2000 174763 287982 175993
rect 2000 172903 287982 174133
rect 2000 169483 287982 172273
rect 2000 167623 287982 168853
rect 2000 165763 287982 166993
rect 2000 163903 287982 165133
rect 2000 160483 287982 163273
rect 2000 158623 287982 159853
rect 2000 156763 287982 157993
rect 2000 154903 287982 156133
rect 2000 151483 287982 154273
rect 2000 149623 287982 150853
rect 2000 147763 287982 148993
rect 2000 145903 287982 147133
rect 2000 142483 287982 145273
rect 2000 140623 287982 141853
rect 2000 138763 287982 139993
rect 2000 136903 287982 138133
rect 2000 133483 287982 136273
rect 2000 131623 287982 132853
rect 2000 129763 287982 130993
rect 2000 127903 287982 129133
rect 2000 124483 287982 127273
rect 2000 122623 287982 123853
rect 2000 120763 287982 121993
rect 2000 118903 287982 120133
rect 2000 115483 287982 118273
rect 2000 113623 287982 114853
rect 2000 111763 287982 112993
rect 2000 109903 287982 111133
rect 2000 106483 287982 109273
rect 2000 104623 287982 105853
rect 2000 102763 287982 103993
rect 2000 100903 287982 102133
rect 2000 97483 287982 100273
rect 2000 95623 287982 96853
rect 2000 93763 287982 94993
rect 2000 91903 287982 93133
rect 2000 88483 287982 91273
rect 2000 86623 287982 87853
rect 2000 84763 287982 85993
rect 2000 82903 287982 84133
rect 2000 79483 287982 82273
rect 2000 77623 287982 78853
rect 2000 75763 287982 76993
rect 2000 73903 287982 75133
rect 2000 70483 287982 73273
rect 2000 68623 287982 69853
rect 2000 66763 287982 67993
rect 2000 64903 287982 66133
rect 2000 61483 287982 64273
rect 2000 59623 287982 60853
rect 2000 57763 287982 58993
rect 2000 55903 287982 57133
rect 2000 52483 287982 55273
rect 2000 50623 287982 51853
rect 2000 48763 287982 49993
rect 2000 46903 287982 48133
rect 2000 43483 287982 46273
rect 2000 41623 287982 42853
rect 2000 39763 287982 40993
rect 2000 37903 287982 39133
rect 2000 34483 287982 37273
rect 2000 32623 287982 33853
rect 2000 30763 287982 31993
rect 2000 28903 287982 30133
rect 2000 25483 287982 28273
rect 2000 23623 287982 24853
rect 2000 21763 287982 22993
rect 2000 19903 287982 21133
rect 2000 16483 287982 19273
rect 2000 14623 287982 15853
rect 2000 12763 287982 13993
rect 2000 10903 287982 12133
rect 2000 7483 287982 10273
rect 2000 5623 287982 6853
rect 2000 3926 287982 4993
<< labels >>
rlabel metal3 s 291760 142638 292480 142758 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 223049 351760 223105 352480 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 190573 351760 190629 352480 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 158143 351760 158199 352480 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 125713 351760 125769 352480 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 93237 351760 93293 352480 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 60807 351760 60863 352480 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 28377 351760 28433 352480 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -480 348610 240 348730 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -480 322498 240 322618 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -480 296454 240 296574 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 291760 169226 292480 169346 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -480 270342 240 270462 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -480 244298 240 244418 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -480 218254 240 218374 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -480 192142 240 192262 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -480 166098 240 166218 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -480 139986 240 140106 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -480 113942 240 114062 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -480 87898 240 88018 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -480 61786 240 61906 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 291760 195814 292480 195934 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 291760 222334 292480 222454 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 291760 248922 292480 249042 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 291760 275510 292480 275630 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 291760 302030 292480 302150 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 291760 328618 292480 328738 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 287909 351760 287965 352480 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 255479 351760 255535 352480 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 291760 3238 292480 3358 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 291760 228998 292480 229118 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 291760 255586 292480 255706 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 291760 282106 292480 282226 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 291760 308694 292480 308814 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 291760 335282 292480 335402 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 279813 351760 279869 352480 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 247383 351760 247439 352480 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 214907 351760 214963 352480 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 182477 351760 182533 352480 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 150047 351760 150103 352480 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 291760 23094 292480 23214 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 117571 351760 117627 352480 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 85141 351760 85197 352480 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 52711 351760 52767 352480 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 20235 351760 20291 352480 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -480 342082 240 342202 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -480 315970 240 316090 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -480 289926 240 290046 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -480 263882 240 264002 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -480 237770 240 237890 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -480 211726 240 211846 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 291760 43018 292480 43138 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -480 185614 240 185734 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -480 159570 240 159690 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -480 133526 240 133646 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -480 107414 240 107534 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -480 81370 240 81490 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -480 55258 240 55378 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -480 35742 240 35862 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -480 16158 240 16278 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 291760 62942 292480 63062 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 291760 82866 292480 82986 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 291760 102790 292480 102910 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 291760 122714 292480 122834 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 291760 149302 292480 149422 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 291760 175890 292480 176010 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 291760 202410 292480 202530 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 291760 16498 292480 16618 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 291760 242258 292480 242378 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 291760 268846 292480 268966 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 291760 295434 292480 295554 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 291760 321954 292480 322074 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 291760 348542 292480 348662 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 263575 351760 263631 352480 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 231145 351760 231201 352480 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 198715 351760 198771 352480 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 166239 351760 166295 352480 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 133809 351760 133865 352480 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 291760 36422 292480 36542 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 101379 351760 101435 352480 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 68903 351760 68959 352480 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 36473 351760 36529 352480 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 4043 351760 4099 352480 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -480 329026 240 329146 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -480 302982 240 303102 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -480 276870 240 276990 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -480 250826 240 250946 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -480 224714 240 224834 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -480 198670 240 198790 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 291760 56346 292480 56466 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -480 172626 240 172746 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -480 146514 240 146634 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -480 120470 240 120590 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -480 94358 240 94478 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -480 68314 240 68434 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -480 42270 240 42390 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -480 22686 240 22806 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -480 3170 240 3290 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 291760 76270 292480 76390 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 291760 96194 292480 96314 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 291760 116118 292480 116238 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 291760 136042 292480 136162 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 291760 162562 292480 162682 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 291760 189150 292480 189270 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 291760 215738 292480 215858 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 291760 9834 292480 9954 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 291760 235662 292480 235782 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 291760 262182 292480 262302 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 291760 288770 292480 288890 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 291760 315358 292480 315478 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 291760 341878 292480 341998 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 271717 351760 271773 352480 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 239241 351760 239297 352480 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 206811 351760 206867 352480 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 174381 351760 174437 352480 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 141905 351760 141961 352480 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 291760 29758 292480 29878 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 109475 351760 109531 352480 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 77045 351760 77101 352480 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 44569 351760 44625 352480 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 12139 351760 12195 352480 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -480 335554 240 335674 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -480 309510 240 309630 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -480 283398 240 283518 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -480 257354 240 257474 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -480 231242 240 231362 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -480 205198 240 205318 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 291760 49682 292480 49802 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -480 179154 240 179274 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -480 153042 240 153162 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -480 126998 240 127118 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -480 100886 240 101006 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -480 74842 240 74962 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -480 48730 240 48850 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -480 29214 240 29334 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -480 9630 240 9750 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 291760 69606 292480 69726 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 291760 89530 292480 89650 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 291760 109454 292480 109574 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 291760 129378 292480 129498 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 291760 155966 292480 156086 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 291760 182486 292480 182606 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 291760 209074 292480 209194 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 62923 -480 62979 240 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 240253 -480 240309 240 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 242001 -480 242057 240 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 243795 -480 243851 240 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 245543 -480 245599 240 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 247337 -480 247393 240 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 249085 -480 249141 240 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 250879 -480 250935 240 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 252673 -480 252729 240 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 254421 -480 254477 240 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 256215 -480 256271 240 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 80633 -480 80689 240 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 257963 -480 258019 240 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 259757 -480 259813 240 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 261505 -480 261561 240 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 263299 -480 263355 240 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 265047 -480 265103 240 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 266841 -480 266897 240 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 268589 -480 268645 240 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 270383 -480 270439 240 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 272177 -480 272233 240 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 273925 -480 273981 240 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 82427 -480 82483 240 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 275719 -480 275775 240 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 277467 -480 277523 240 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 279261 -480 279317 240 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 281009 -480 281065 240 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 282803 -480 282859 240 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 284551 -480 284607 240 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 286345 -480 286401 240 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 288139 -480 288195 240 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 84175 -480 84231 240 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 85969 -480 86025 240 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 87717 -480 87773 240 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 89511 -480 89567 240 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 91259 -480 91315 240 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 93053 -480 93109 240 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 94847 -480 94903 240 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 96595 -480 96651 240 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 64671 -480 64727 240 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 98389 -480 98445 240 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 100137 -480 100193 240 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 101931 -480 101987 240 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 103679 -480 103735 240 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 105473 -480 105529 240 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 107221 -480 107277 240 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 109015 -480 109071 240 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 110763 -480 110819 240 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 112557 -480 112613 240 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 114351 -480 114407 240 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 66465 -480 66521 240 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 116099 -480 116155 240 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 117893 -480 117949 240 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 119641 -480 119697 240 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 121435 -480 121491 240 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 123183 -480 123239 240 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 124977 -480 125033 240 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 126725 -480 126781 240 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 128519 -480 128575 240 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 130313 -480 130369 240 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 132061 -480 132117 240 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 68213 -480 68269 240 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 133855 -480 133911 240 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 135603 -480 135659 240 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 137397 -480 137453 240 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 139145 -480 139201 240 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 140939 -480 140995 240 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 142687 -480 142743 240 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 144481 -480 144537 240 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 146275 -480 146331 240 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 148023 -480 148079 240 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 149817 -480 149873 240 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 70007 -480 70063 240 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 151565 -480 151621 240 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 153359 -480 153415 240 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 155107 -480 155163 240 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 156901 -480 156957 240 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 158649 -480 158705 240 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 160443 -480 160499 240 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 162191 -480 162247 240 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 163985 -480 164041 240 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 165779 -480 165835 240 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 167527 -480 167583 240 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 71755 -480 71811 240 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 169321 -480 169377 240 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 171069 -480 171125 240 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 172863 -480 172919 240 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 174611 -480 174667 240 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 176405 -480 176461 240 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 178153 -480 178209 240 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 179947 -480 180003 240 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 181741 -480 181797 240 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 183489 -480 183545 240 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 185283 -480 185339 240 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 73549 -480 73605 240 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 187031 -480 187087 240 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 188825 -480 188881 240 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 190573 -480 190629 240 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 192367 -480 192423 240 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 194115 -480 194171 240 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 195909 -480 195965 240 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 197657 -480 197713 240 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 199451 -480 199507 240 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 201245 -480 201301 240 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 202993 -480 203049 240 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 75297 -480 75353 240 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 204787 -480 204843 240 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 206535 -480 206591 240 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 208329 -480 208385 240 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 210077 -480 210133 240 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 211871 -480 211927 240 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 213619 -480 213675 240 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 215413 -480 215469 240 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 217207 -480 217263 240 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 218955 -480 219011 240 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 220749 -480 220805 240 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 77091 -480 77147 240 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 222497 -480 222553 240 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 224291 -480 224347 240 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 226039 -480 226095 240 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 227833 -480 227889 240 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 229581 -480 229637 240 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 231375 -480 231431 240 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 233123 -480 233179 240 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 234917 -480 234973 240 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 236711 -480 236767 240 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 238459 -480 238515 240 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 78885 -480 78941 240 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 63475 -480 63531 240 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 240851 -480 240907 240 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 242599 -480 242655 240 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 244393 -480 244449 240 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 246141 -480 246197 240 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 247935 -480 247991 240 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 249683 -480 249739 240 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 251477 -480 251533 240 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 253225 -480 253281 240 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 255019 -480 255075 240 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 256767 -480 256823 240 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 81231 -480 81287 240 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 258561 -480 258617 240 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 260355 -480 260411 240 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 262103 -480 262159 240 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 263897 -480 263953 240 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 265645 -480 265701 240 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 267439 -480 267495 240 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 269187 -480 269243 240 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 270981 -480 271037 240 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 272729 -480 272785 240 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 274523 -480 274579 240 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 83025 -480 83081 240 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 276317 -480 276373 240 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 278065 -480 278121 240 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 279859 -480 279915 240 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 281607 -480 281663 240 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 283401 -480 283457 240 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 285149 -480 285205 240 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 286943 -480 286999 240 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 288691 -480 288747 240 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 84773 -480 84829 240 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 86567 -480 86623 240 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 88315 -480 88371 240 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 90109 -480 90165 240 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 91857 -480 91913 240 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 93651 -480 93707 240 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 95399 -480 95455 240 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 97193 -480 97249 240 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 65269 -480 65325 240 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 98941 -480 98997 240 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 100735 -480 100791 240 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 102529 -480 102585 240 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 104277 -480 104333 240 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 106071 -480 106127 240 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 107819 -480 107875 240 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 109613 -480 109669 240 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 111361 -480 111417 240 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 113155 -480 113211 240 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 114903 -480 114959 240 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 67063 -480 67119 240 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 116697 -480 116753 240 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 118491 -480 118547 240 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 120239 -480 120295 240 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 122033 -480 122089 240 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 123781 -480 123837 240 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 125575 -480 125631 240 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 127323 -480 127379 240 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 129117 -480 129173 240 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 130865 -480 130921 240 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 132659 -480 132715 240 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 68811 -480 68867 240 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 134407 -480 134463 240 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 136201 -480 136257 240 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 137995 -480 138051 240 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 139743 -480 139799 240 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 141537 -480 141593 240 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 143285 -480 143341 240 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 145079 -480 145135 240 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 146827 -480 146883 240 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 148621 -480 148677 240 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 150369 -480 150425 240 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 70605 -480 70661 240 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 152163 -480 152219 240 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 153957 -480 154013 240 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 155705 -480 155761 240 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 157499 -480 157555 240 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 159247 -480 159303 240 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 161041 -480 161097 240 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 162789 -480 162845 240 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 164583 -480 164639 240 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 166331 -480 166387 240 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 168125 -480 168181 240 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 72353 -480 72409 240 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 169919 -480 169975 240 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 171667 -480 171723 240 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 173461 -480 173517 240 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 175209 -480 175265 240 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 177003 -480 177059 240 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 178751 -480 178807 240 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 180545 -480 180601 240 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 182293 -480 182349 240 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 184087 -480 184143 240 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 185835 -480 185891 240 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 74147 -480 74203 240 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 187629 -480 187685 240 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 189423 -480 189479 240 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 191171 -480 191227 240 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 192965 -480 193021 240 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 194713 -480 194769 240 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 196507 -480 196563 240 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 198255 -480 198311 240 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 200049 -480 200105 240 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 201797 -480 201853 240 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 203591 -480 203647 240 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 75895 -480 75951 240 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 205385 -480 205441 240 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 207133 -480 207189 240 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 208927 -480 208983 240 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 210675 -480 210731 240 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 212469 -480 212525 240 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 214217 -480 214273 240 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 216011 -480 216067 240 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 217759 -480 217815 240 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 219553 -480 219609 240 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 221301 -480 221357 240 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 77689 -480 77745 240 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 223095 -480 223151 240 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 224889 -480 224945 240 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 226637 -480 226693 240 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 228431 -480 228487 240 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 230179 -480 230235 240 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 231973 -480 232029 240 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 233721 -480 233777 240 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 235515 -480 235571 240 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 237263 -480 237319 240 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 239057 -480 239113 240 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 79437 -480 79493 240 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 64073 -480 64129 240 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 241403 -480 241459 240 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 243197 -480 243253 240 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 244945 -480 245001 240 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 246739 -480 246795 240 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 248533 -480 248589 240 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 250281 -480 250337 240 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 252075 -480 252131 240 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 253823 -480 253879 240 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 255617 -480 255673 240 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 257365 -480 257421 240 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 81829 -480 81885 240 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 259159 -480 259215 240 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 260907 -480 260963 240 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 262701 -480 262757 240 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 264495 -480 264551 240 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 266243 -480 266299 240 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 268037 -480 268093 240 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 269785 -480 269841 240 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 271579 -480 271635 240 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 273327 -480 273383 240 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 275121 -480 275177 240 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 83577 -480 83633 240 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 276869 -480 276925 240 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 278663 -480 278719 240 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 280411 -480 280467 240 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 282205 -480 282261 240 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 283999 -480 284055 240 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 285747 -480 285803 240 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 287541 -480 287597 240 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 289289 -480 289345 240 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 85371 -480 85427 240 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 87119 -480 87175 240 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 88913 -480 88969 240 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 90707 -480 90763 240 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 92455 -480 92511 240 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 94249 -480 94305 240 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 95997 -480 96053 240 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 97791 -480 97847 240 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 65867 -480 65923 240 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 99539 -480 99595 240 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 101333 -480 101389 240 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 103081 -480 103137 240 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 104875 -480 104931 240 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 106669 -480 106725 240 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 108417 -480 108473 240 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 110211 -480 110267 240 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 111959 -480 112015 240 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 113753 -480 113809 240 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 115501 -480 115557 240 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 67615 -480 67671 240 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 117295 -480 117351 240 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 119043 -480 119099 240 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 120837 -480 120893 240 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 122585 -480 122641 240 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 124379 -480 124435 240 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 126173 -480 126229 240 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 127921 -480 127977 240 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 129715 -480 129771 240 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 131463 -480 131519 240 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 133257 -480 133313 240 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 69409 -480 69465 240 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 135005 -480 135061 240 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 136799 -480 136855 240 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 138547 -480 138603 240 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 140341 -480 140397 240 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 142135 -480 142191 240 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 143883 -480 143939 240 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 145677 -480 145733 240 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 147425 -480 147481 240 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 149219 -480 149275 240 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 150967 -480 151023 240 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 71203 -480 71259 240 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 152761 -480 152817 240 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 154509 -480 154565 240 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 156303 -480 156359 240 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 158097 -480 158153 240 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 159845 -480 159901 240 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 161639 -480 161695 240 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 163387 -480 163443 240 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 165181 -480 165237 240 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 166929 -480 166985 240 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 168723 -480 168779 240 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 72951 -480 73007 240 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 170471 -480 170527 240 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 172265 -480 172321 240 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 174013 -480 174069 240 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 175807 -480 175863 240 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 177601 -480 177657 240 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 179349 -480 179405 240 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 181143 -480 181199 240 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 182891 -480 182947 240 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 184685 -480 184741 240 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 186433 -480 186489 240 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 74745 -480 74801 240 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 188227 -480 188283 240 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 189975 -480 190031 240 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 191769 -480 191825 240 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 193563 -480 193619 240 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 195311 -480 195367 240 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 197105 -480 197161 240 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 198853 -480 198909 240 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 200647 -480 200703 240 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 202395 -480 202451 240 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 204189 -480 204245 240 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 76493 -480 76549 240 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 205937 -480 205993 240 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 207731 -480 207787 240 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 209479 -480 209535 240 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 211273 -480 211329 240 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 213067 -480 213123 240 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 214815 -480 214871 240 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 216609 -480 216665 240 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 218357 -480 218413 240 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 220151 -480 220207 240 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 221899 -480 221955 240 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 78287 -480 78343 240 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 223693 -480 223749 240 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 225441 -480 225497 240 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 227235 -480 227291 240 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 229029 -480 229085 240 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 230777 -480 230833 240 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 232571 -480 232627 240 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 234319 -480 234375 240 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 236113 -480 236169 240 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 237861 -480 237917 240 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 239655 -480 239711 240 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 80035 -480 80091 240 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 289887 -480 289943 240 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 290485 -480 290541 240 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 291083 -480 291139 240 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 291681 -480 291737 240 8 user_irq[2]
port 531 nsew signal output
rlabel metal5 s -1003 -467 292965 -157 8 vccd1
port 532 nsew power input
rlabel metal5 s -1483 1433 293445 1743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 19433 293445 19743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 37433 293445 37743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 55433 293445 55743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 73433 293445 73743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 91433 293445 91743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 109433 293445 109743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 127433 293445 127743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 145433 293445 145743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 163433 293445 163743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 181433 293445 181743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 199433 293445 199743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 217433 293445 217743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 235433 293445 235743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 253433 293445 253743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 271433 293445 271743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 289433 293445 289743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 307433 293445 307743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 325433 293445 325743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1483 343433 293445 343743 6 vccd1
port 532 nsew power input
rlabel metal5 s -1003 352125 292965 352435 6 vccd1
port 532 nsew power input
rlabel metal4 s 897 -947 1207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 18897 -947 19207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 36897 -947 37207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 54897 -947 55207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 72897 -947 73207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 90897 -947 91207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 108897 -947 109207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 126897 -947 127207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 144897 -947 145207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 162897 -947 163207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 180897 -947 181207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 198897 -947 199207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 216897 -947 217207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 234897 -947 235207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 252897 -947 253207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 270897 -947 271207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s 288897 -947 289207 1000 6 vccd1
port 532 nsew power input
rlabel metal4 s -1003 -467 -693 352435 4 vccd1
port 532 nsew power input
rlabel metal4 s 292655 -467 292965 352435 6 vccd1
port 532 nsew power input
rlabel metal4 s 897 350004 1207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 18897 350004 19207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 36897 350004 37207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 54897 350004 55207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 72897 350004 73207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 90897 350004 91207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 108897 350004 109207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 126897 350004 127207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 144897 350004 145207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 162897 350004 163207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 180897 350004 181207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 198897 350004 199207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 216897 350004 217207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 234897 350004 235207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 252897 350004 253207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 270897 350004 271207 352915 6 vccd1
port 532 nsew power input
rlabel metal4 s 288897 350004 289207 352915 6 vccd1
port 532 nsew power input
rlabel metal5 s -1963 -1427 293925 -1117 8 vccd2
port 533 nsew power input
rlabel metal5 s -2443 3293 294405 3603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 21293 294405 21603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 39293 294405 39603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 57293 294405 57603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 75293 294405 75603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 93293 294405 93603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 111293 294405 111603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 129293 294405 129603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 147293 294405 147603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 165293 294405 165603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 183293 294405 183603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 201293 294405 201603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 219293 294405 219603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 237293 294405 237603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 255293 294405 255603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 273293 294405 273603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 291293 294405 291603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 309293 294405 309603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 327293 294405 327603 6 vccd2
port 533 nsew power input
rlabel metal5 s -2443 345293 294405 345603 6 vccd2
port 533 nsew power input
rlabel metal5 s -1963 353085 293925 353395 6 vccd2
port 533 nsew power input
rlabel metal4 s 2757 -1907 3067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s 20757 -1907 21067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s 38757 -1907 39067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s 56757 -1907 57067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s 74757 -1907 75067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s 92757 -1907 93067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s 110757 -1907 111067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s 128757 -1907 129067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s 146757 -1907 147067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s 164757 -1907 165067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s 182757 -1907 183067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s 200757 -1907 201067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s 218757 -1907 219067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s 236757 -1907 237067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s 254757 -1907 255067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s 272757 -1907 273067 1000 8 vccd2
port 533 nsew power input
rlabel metal4 s -1963 -1427 -1653 353395 4 vccd2
port 533 nsew power input
rlabel metal4 s 293615 -1427 293925 353395 6 vccd2
port 533 nsew power input
rlabel metal4 s 2757 350004 3067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 20757 350004 21067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 38757 350004 39067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 56757 350004 57067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 74757 350004 75067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 92757 350004 93067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 110757 350004 111067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 128757 350004 129067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 146757 350004 147067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 164757 350004 165067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 182757 350004 183067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 200757 350004 201067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 218757 350004 219067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 236757 350004 237067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 254757 350004 255067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 272757 350004 273067 353875 6 vccd2
port 533 nsew power input
rlabel metal4 s 290757 -1907 291067 353875 6 vccd2
port 533 nsew power input
rlabel metal5 s -2923 -2387 294885 -2077 8 vdda1
port 534 nsew power input
rlabel metal5 s -3403 5153 295365 5463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 23153 295365 23463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 41153 295365 41463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 59153 295365 59463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 77153 295365 77463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 95153 295365 95463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 113153 295365 113463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 131153 295365 131463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 149153 295365 149463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 167153 295365 167463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 185153 295365 185463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 203153 295365 203463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 221153 295365 221463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 239153 295365 239463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 257153 295365 257463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 275153 295365 275463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 293153 295365 293463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 311153 295365 311463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 329153 295365 329463 6 vdda1
port 534 nsew power input
rlabel metal5 s -3403 347153 295365 347463 6 vdda1
port 534 nsew power input
rlabel metal5 s -2923 354045 294885 354355 6 vdda1
port 534 nsew power input
rlabel metal4 s 4617 -2867 4927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s 22617 -2867 22927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s 40617 -2867 40927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s 58617 -2867 58927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s 76617 -2867 76927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s 94617 -2867 94927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s 112617 -2867 112927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s 130617 -2867 130927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s 148617 -2867 148927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s 166617 -2867 166927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s 184617 -2867 184927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s 202617 -2867 202927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s 220617 -2867 220927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s 238617 -2867 238927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s 256617 -2867 256927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s 274617 -2867 274927 1000 8 vdda1
port 534 nsew power input
rlabel metal4 s -2923 -2387 -2613 354355 4 vdda1
port 534 nsew power input
rlabel metal4 s 294575 -2387 294885 354355 6 vdda1
port 534 nsew power input
rlabel metal4 s 4617 350004 4927 354835 6 vdda1
port 534 nsew power input
rlabel metal4 s 22617 350004 22927 354835 6 vdda1
port 534 nsew power input
rlabel metal4 s 40617 350004 40927 354835 6 vdda1
port 534 nsew power input
rlabel metal4 s 58617 350004 58927 354835 6 vdda1
port 534 nsew power input
rlabel metal4 s 76617 350004 76927 354835 6 vdda1
port 534 nsew power input
rlabel metal4 s 94617 350004 94927 354835 6 vdda1
port 534 nsew power input
rlabel metal4 s 112617 350004 112927 354835 6 vdda1
port 534 nsew power input
rlabel metal4 s 130617 350004 130927 354835 6 vdda1
port 534 nsew power input
rlabel metal4 s 148617 350004 148927 354835 6 vdda1
port 534 nsew power input
rlabel metal4 s 166617 350004 166927 354835 6 vdda1
port 534 nsew power input
rlabel metal4 s 184617 350004 184927 354835 6 vdda1
port 534 nsew power input
rlabel metal4 s 202617 350004 202927 354835 6 vdda1
port 534 nsew power input
rlabel metal4 s 220617 350004 220927 354835 6 vdda1
port 534 nsew power input
rlabel metal4 s 238617 350004 238927 354835 6 vdda1
port 534 nsew power input
rlabel metal4 s 256617 350004 256927 354835 6 vdda1
port 534 nsew power input
rlabel metal4 s 274617 350004 274927 354835 6 vdda1
port 534 nsew power input
rlabel metal5 s -3883 -3347 295845 -3037 8 vdda2
port 535 nsew power input
rlabel metal5 s -4363 7013 296325 7323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 25013 296325 25323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 43013 296325 43323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 61013 296325 61323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 79013 296325 79323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 97013 296325 97323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 115013 296325 115323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 133013 296325 133323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 151013 296325 151323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 169013 296325 169323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 187013 296325 187323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 205013 296325 205323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 223013 296325 223323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 241013 296325 241323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 259013 296325 259323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 277013 296325 277323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 295013 296325 295323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 313013 296325 313323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 331013 296325 331323 6 vdda2
port 535 nsew power input
rlabel metal5 s -4363 349013 296325 349323 6 vdda2
port 535 nsew power input
rlabel metal5 s -3883 355005 295845 355315 6 vdda2
port 535 nsew power input
rlabel metal4 s 6477 -3827 6787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s 24477 -3827 24787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s 42477 -3827 42787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s 60477 -3827 60787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s 78477 -3827 78787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s 96477 -3827 96787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s 114477 -3827 114787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s 132477 -3827 132787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s 150477 -3827 150787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s 168477 -3827 168787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s 186477 -3827 186787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s 204477 -3827 204787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s 222477 -3827 222787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s 240477 -3827 240787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s 258477 -3827 258787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s 276477 -3827 276787 1000 8 vdda2
port 535 nsew power input
rlabel metal4 s -3883 -3347 -3573 355315 4 vdda2
port 535 nsew power input
rlabel metal4 s 295535 -3347 295845 355315 6 vdda2
port 535 nsew power input
rlabel metal4 s 6477 350004 6787 355795 6 vdda2
port 535 nsew power input
rlabel metal4 s 24477 350004 24787 355795 6 vdda2
port 535 nsew power input
rlabel metal4 s 42477 350004 42787 355795 6 vdda2
port 535 nsew power input
rlabel metal4 s 60477 350004 60787 355795 6 vdda2
port 535 nsew power input
rlabel metal4 s 78477 350004 78787 355795 6 vdda2
port 535 nsew power input
rlabel metal4 s 96477 350004 96787 355795 6 vdda2
port 535 nsew power input
rlabel metal4 s 114477 350004 114787 355795 6 vdda2
port 535 nsew power input
rlabel metal4 s 132477 350004 132787 355795 6 vdda2
port 535 nsew power input
rlabel metal4 s 150477 350004 150787 355795 6 vdda2
port 535 nsew power input
rlabel metal4 s 168477 350004 168787 355795 6 vdda2
port 535 nsew power input
rlabel metal4 s 186477 350004 186787 355795 6 vdda2
port 535 nsew power input
rlabel metal4 s 204477 350004 204787 355795 6 vdda2
port 535 nsew power input
rlabel metal4 s 222477 350004 222787 355795 6 vdda2
port 535 nsew power input
rlabel metal4 s 240477 350004 240787 355795 6 vdda2
port 535 nsew power input
rlabel metal4 s 258477 350004 258787 355795 6 vdda2
port 535 nsew power input
rlabel metal4 s 276477 350004 276787 355795 6 vdda2
port 535 nsew power input
rlabel metal5 s -3403 -2867 295365 -2557 8 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 14153 295365 14463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 32153 295365 32463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 50153 295365 50463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 68153 295365 68463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 86153 295365 86463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 104153 295365 104463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 122153 295365 122463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 140153 295365 140463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 158153 295365 158463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 176153 295365 176463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 194153 295365 194463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 212153 295365 212463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 230153 295365 230463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 248153 295365 248463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 266153 295365 266463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 284153 295365 284463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 302153 295365 302463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 320153 295365 320463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 338153 295365 338463 6 vssa1
port 536 nsew ground input
rlabel metal5 s -3403 354525 295365 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 13617 -2867 13927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 31617 -2867 31927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 49617 -2867 49927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 67617 -2867 67927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 85617 -2867 85927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 103617 -2867 103927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 121617 -2867 121927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 139617 -2867 139927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 157617 -2867 157927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 175617 -2867 175927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 193617 -2867 193927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 211617 -2867 211927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 229617 -2867 229927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 247617 -2867 247927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 265617 -2867 265927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 283617 -2867 283927 1000 8 vssa1
port 536 nsew ground input
rlabel metal4 s -3403 -2867 -3093 354835 4 vssa1
port 536 nsew ground input
rlabel metal4 s 13617 350004 13927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 31617 350004 31927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 49617 350004 49927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 67617 350004 67927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 85617 350004 85927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 103617 350004 103927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 121617 350004 121927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 139617 350004 139927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 157617 350004 157927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 175617 350004 175927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 193617 350004 193927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 211617 350004 211927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 229617 350004 229927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 247617 350004 247927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 265617 350004 265927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 283617 350004 283927 354835 6 vssa1
port 536 nsew ground input
rlabel metal4 s 295055 -2867 295365 354835 6 vssa1
port 536 nsew ground input
rlabel metal5 s -4363 -3827 296325 -3517 8 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 16013 296325 16323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 34013 296325 34323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 52013 296325 52323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 70013 296325 70323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 88013 296325 88323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 106013 296325 106323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 124013 296325 124323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 142013 296325 142323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 160013 296325 160323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 178013 296325 178323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 196013 296325 196323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 214013 296325 214323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 232013 296325 232323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 250013 296325 250323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 268013 296325 268323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 286013 296325 286323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 304013 296325 304323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 322013 296325 322323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 340013 296325 340323 6 vssa2
port 537 nsew ground input
rlabel metal5 s -4363 355485 296325 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 15477 -3827 15787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 33477 -3827 33787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 51477 -3827 51787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 69477 -3827 69787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 87477 -3827 87787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 105477 -3827 105787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 123477 -3827 123787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 141477 -3827 141787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 159477 -3827 159787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 177477 -3827 177787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 195477 -3827 195787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 213477 -3827 213787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 231477 -3827 231787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 249477 -3827 249787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 267477 -3827 267787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 285477 -3827 285787 1000 8 vssa2
port 537 nsew ground input
rlabel metal4 s -4363 -3827 -4053 355795 4 vssa2
port 537 nsew ground input
rlabel metal4 s 15477 350004 15787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 33477 350004 33787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 51477 350004 51787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 69477 350004 69787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 87477 350004 87787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 105477 350004 105787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 123477 350004 123787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 141477 350004 141787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 159477 350004 159787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 177477 350004 177787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 195477 350004 195787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 213477 350004 213787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 231477 350004 231787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 249477 350004 249787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 267477 350004 267787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 285477 350004 285787 355795 6 vssa2
port 537 nsew ground input
rlabel metal4 s 296015 -3827 296325 355795 6 vssa2
port 537 nsew ground input
rlabel metal5 s -1483 -947 293445 -637 8 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 10433 293445 10743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 28433 293445 28743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 46433 293445 46743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 64433 293445 64743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 82433 293445 82743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 100433 293445 100743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 118433 293445 118743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 136433 293445 136743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 154433 293445 154743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 172433 293445 172743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 190433 293445 190743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 208433 293445 208743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 226433 293445 226743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 244433 293445 244743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 262433 293445 262743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 280433 293445 280743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 298433 293445 298743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 316433 293445 316743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 334433 293445 334743 6 vssd1
port 538 nsew ground input
rlabel metal5 s -1483 352605 293445 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 9897 -947 10207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 27897 -947 28207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 45897 -947 46207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 63897 -947 64207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 81897 -947 82207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 99897 -947 100207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 117897 -947 118207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 135897 -947 136207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 153897 -947 154207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 171897 -947 172207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 189897 -947 190207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 207897 -947 208207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 225897 -947 226207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 243897 -947 244207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 261897 -947 262207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 279897 -947 280207 1000 6 vssd1
port 538 nsew ground input
rlabel metal4 s -1483 -947 -1173 352915 4 vssd1
port 538 nsew ground input
rlabel metal4 s 9897 350004 10207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 27897 350004 28207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 45897 350004 46207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 63897 350004 64207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 81897 350004 82207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 99897 350004 100207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 117897 350004 118207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 135897 350004 136207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 153897 350004 154207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 171897 350004 172207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 189897 350004 190207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 207897 350004 208207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 225897 350004 226207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 243897 350004 244207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 261897 350004 262207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 279897 350004 280207 352915 6 vssd1
port 538 nsew ground input
rlabel metal4 s 293135 -947 293445 352915 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2443 -1907 294405 -1597 8 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 12293 294405 12603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 30293 294405 30603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 48293 294405 48603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 66293 294405 66603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 84293 294405 84603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 102293 294405 102603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 120293 294405 120603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 138293 294405 138603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 156293 294405 156603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 174293 294405 174603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 192293 294405 192603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 210293 294405 210603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 228293 294405 228603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 246293 294405 246603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 264293 294405 264603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 282293 294405 282603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 300293 294405 300603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 318293 294405 318603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 336293 294405 336603 6 vssd2
port 539 nsew ground input
rlabel metal5 s -2443 353565 294405 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 11757 -1907 12067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s 29757 -1907 30067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s 47757 -1907 48067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s 65757 -1907 66067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s 83757 -1907 84067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s 101757 -1907 102067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s 119757 -1907 120067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s 137757 -1907 138067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s 155757 -1907 156067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s 173757 -1907 174067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s 191757 -1907 192067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s 209757 -1907 210067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s 227757 -1907 228067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s 245757 -1907 246067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s 263757 -1907 264067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s 281757 -1907 282067 1000 8 vssd2
port 539 nsew ground input
rlabel metal4 s -2443 -1907 -2133 353875 4 vssd2
port 539 nsew ground input
rlabel metal4 s 11757 350004 12067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 29757 350004 30067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 47757 350004 48067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 65757 350004 66067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 83757 350004 84067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 101757 350004 102067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 119757 350004 120067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 137757 350004 138067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 155757 350004 156067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 173757 350004 174067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 191757 350004 192067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 209757 350004 210067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 227757 350004 228067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 245757 350004 246067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 263757 350004 264067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 281757 350004 282067 353875 6 vssd2
port 539 nsew ground input
rlabel metal4 s 294095 -1907 294405 353875 6 vssd2
port 539 nsew ground input
rlabel metal2 s 271 -480 327 240 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 823 -480 879 240 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 1421 -480 1477 240 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 3813 -480 3869 240 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 23915 -480 23971 240 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 25663 -480 25719 240 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 27457 -480 27513 240 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 29205 -480 29261 240 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 30999 -480 31055 240 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 32747 -480 32803 240 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 34541 -480 34597 240 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 36289 -480 36345 240 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 38083 -480 38139 240 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 39831 -480 39887 240 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 6159 -480 6215 240 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 41625 -480 41681 240 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 43419 -480 43475 240 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 45167 -480 45223 240 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 46961 -480 47017 240 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 48709 -480 48765 240 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 50503 -480 50559 240 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 52251 -480 52307 240 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 54045 -480 54101 240 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 55793 -480 55849 240 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 57587 -480 57643 240 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 8505 -480 8561 240 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 59381 -480 59437 240 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 61129 -480 61185 240 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 10897 -480 10953 240 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 13243 -480 13299 240 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 15037 -480 15093 240 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 16785 -480 16841 240 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 18579 -480 18635 240 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 20327 -480 20383 240 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 22121 -480 22177 240 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 2019 -480 2075 240 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 4365 -480 4421 240 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 24467 -480 24523 240 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 26261 -480 26317 240 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 28009 -480 28065 240 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 29803 -480 29859 240 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 31597 -480 31653 240 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 33345 -480 33401 240 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 35139 -480 35195 240 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 36887 -480 36943 240 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 38681 -480 38737 240 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 40429 -480 40485 240 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 6757 -480 6813 240 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 42223 -480 42279 240 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 43971 -480 44027 240 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 45765 -480 45821 240 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 47559 -480 47615 240 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 49307 -480 49363 240 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 51101 -480 51157 240 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 52849 -480 52905 240 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 54643 -480 54699 240 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 56391 -480 56447 240 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 58185 -480 58241 240 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 9103 -480 9159 240 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 59933 -480 59989 240 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 61727 -480 61783 240 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 11495 -480 11551 240 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 13841 -480 13897 240 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 15635 -480 15691 240 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 17383 -480 17439 240 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 19177 -480 19233 240 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 20925 -480 20981 240 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 22719 -480 22775 240 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 4963 -480 5019 240 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 25065 -480 25121 240 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 26859 -480 26915 240 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 28607 -480 28663 240 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 30401 -480 30457 240 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 32149 -480 32205 240 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 33943 -480 33999 240 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 35737 -480 35793 240 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 37485 -480 37541 240 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 39279 -480 39335 240 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 41027 -480 41083 240 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 7355 -480 7411 240 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 42821 -480 42877 240 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 44569 -480 44625 240 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 46363 -480 46419 240 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 48111 -480 48167 240 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 49905 -480 49961 240 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 51653 -480 51709 240 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 53447 -480 53503 240 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 55241 -480 55297 240 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 56989 -480 57045 240 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 58783 -480 58839 240 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 9701 -480 9757 240 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 60531 -480 60587 240 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 62325 -480 62381 240 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 12093 -480 12149 240 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 14439 -480 14495 240 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 16187 -480 16243 240 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 17981 -480 18037 240 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 19775 -480 19831 240 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 21523 -480 21579 240 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 23317 -480 23373 240 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 5561 -480 5617 240 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 7953 -480 8009 240 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 10299 -480 10355 240 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 12645 -480 12701 240 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 2617 -480 2673 240 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 3215 -480 3271 240 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 292000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 616145150
string GDS_FILE /farmshare/scratch/users/yuchenm/kairos-caravel/openlane/user_project_wrapper/runs/user_project_wrapper/results/finishing/user_project_wrapper.magic.gds
string GDS_START 615111302
<< end >>

